magic
tech sky130A
magscale 1 2
timestamp 1723380300
<< pwell >>
rect -5685 -1210 5685 1210
<< nmos >>
rect -5489 -1000 -5369 1000
rect -5311 -1000 -5191 1000
rect -5133 -1000 -5013 1000
rect -4955 -1000 -4835 1000
rect -4777 -1000 -4657 1000
rect -4599 -1000 -4479 1000
rect -4421 -1000 -4301 1000
rect -4243 -1000 -4123 1000
rect -4065 -1000 -3945 1000
rect -3887 -1000 -3767 1000
rect -3709 -1000 -3589 1000
rect -3531 -1000 -3411 1000
rect -3353 -1000 -3233 1000
rect -3175 -1000 -3055 1000
rect -2997 -1000 -2877 1000
rect -2819 -1000 -2699 1000
rect -2641 -1000 -2521 1000
rect -2463 -1000 -2343 1000
rect -2285 -1000 -2165 1000
rect -2107 -1000 -1987 1000
rect -1929 -1000 -1809 1000
rect -1751 -1000 -1631 1000
rect -1573 -1000 -1453 1000
rect -1395 -1000 -1275 1000
rect -1217 -1000 -1097 1000
rect -1039 -1000 -919 1000
rect -861 -1000 -741 1000
rect -683 -1000 -563 1000
rect -505 -1000 -385 1000
rect -327 -1000 -207 1000
rect -149 -1000 -29 1000
rect 29 -1000 149 1000
rect 207 -1000 327 1000
rect 385 -1000 505 1000
rect 563 -1000 683 1000
rect 741 -1000 861 1000
rect 919 -1000 1039 1000
rect 1097 -1000 1217 1000
rect 1275 -1000 1395 1000
rect 1453 -1000 1573 1000
rect 1631 -1000 1751 1000
rect 1809 -1000 1929 1000
rect 1987 -1000 2107 1000
rect 2165 -1000 2285 1000
rect 2343 -1000 2463 1000
rect 2521 -1000 2641 1000
rect 2699 -1000 2819 1000
rect 2877 -1000 2997 1000
rect 3055 -1000 3175 1000
rect 3233 -1000 3353 1000
rect 3411 -1000 3531 1000
rect 3589 -1000 3709 1000
rect 3767 -1000 3887 1000
rect 3945 -1000 4065 1000
rect 4123 -1000 4243 1000
rect 4301 -1000 4421 1000
rect 4479 -1000 4599 1000
rect 4657 -1000 4777 1000
rect 4835 -1000 4955 1000
rect 5013 -1000 5133 1000
rect 5191 -1000 5311 1000
rect 5369 -1000 5489 1000
<< ndiff >>
rect -5547 988 -5489 1000
rect -5547 -988 -5535 988
rect -5501 -988 -5489 988
rect -5547 -1000 -5489 -988
rect -5369 988 -5311 1000
rect -5369 -988 -5357 988
rect -5323 -988 -5311 988
rect -5369 -1000 -5311 -988
rect -5191 988 -5133 1000
rect -5191 -988 -5179 988
rect -5145 -988 -5133 988
rect -5191 -1000 -5133 -988
rect -5013 988 -4955 1000
rect -5013 -988 -5001 988
rect -4967 -988 -4955 988
rect -5013 -1000 -4955 -988
rect -4835 988 -4777 1000
rect -4835 -988 -4823 988
rect -4789 -988 -4777 988
rect -4835 -1000 -4777 -988
rect -4657 988 -4599 1000
rect -4657 -988 -4645 988
rect -4611 -988 -4599 988
rect -4657 -1000 -4599 -988
rect -4479 988 -4421 1000
rect -4479 -988 -4467 988
rect -4433 -988 -4421 988
rect -4479 -1000 -4421 -988
rect -4301 988 -4243 1000
rect -4301 -988 -4289 988
rect -4255 -988 -4243 988
rect -4301 -1000 -4243 -988
rect -4123 988 -4065 1000
rect -4123 -988 -4111 988
rect -4077 -988 -4065 988
rect -4123 -1000 -4065 -988
rect -3945 988 -3887 1000
rect -3945 -988 -3933 988
rect -3899 -988 -3887 988
rect -3945 -1000 -3887 -988
rect -3767 988 -3709 1000
rect -3767 -988 -3755 988
rect -3721 -988 -3709 988
rect -3767 -1000 -3709 -988
rect -3589 988 -3531 1000
rect -3589 -988 -3577 988
rect -3543 -988 -3531 988
rect -3589 -1000 -3531 -988
rect -3411 988 -3353 1000
rect -3411 -988 -3399 988
rect -3365 -988 -3353 988
rect -3411 -1000 -3353 -988
rect -3233 988 -3175 1000
rect -3233 -988 -3221 988
rect -3187 -988 -3175 988
rect -3233 -1000 -3175 -988
rect -3055 988 -2997 1000
rect -3055 -988 -3043 988
rect -3009 -988 -2997 988
rect -3055 -1000 -2997 -988
rect -2877 988 -2819 1000
rect -2877 -988 -2865 988
rect -2831 -988 -2819 988
rect -2877 -1000 -2819 -988
rect -2699 988 -2641 1000
rect -2699 -988 -2687 988
rect -2653 -988 -2641 988
rect -2699 -1000 -2641 -988
rect -2521 988 -2463 1000
rect -2521 -988 -2509 988
rect -2475 -988 -2463 988
rect -2521 -1000 -2463 -988
rect -2343 988 -2285 1000
rect -2343 -988 -2331 988
rect -2297 -988 -2285 988
rect -2343 -1000 -2285 -988
rect -2165 988 -2107 1000
rect -2165 -988 -2153 988
rect -2119 -988 -2107 988
rect -2165 -1000 -2107 -988
rect -1987 988 -1929 1000
rect -1987 -988 -1975 988
rect -1941 -988 -1929 988
rect -1987 -1000 -1929 -988
rect -1809 988 -1751 1000
rect -1809 -988 -1797 988
rect -1763 -988 -1751 988
rect -1809 -1000 -1751 -988
rect -1631 988 -1573 1000
rect -1631 -988 -1619 988
rect -1585 -988 -1573 988
rect -1631 -1000 -1573 -988
rect -1453 988 -1395 1000
rect -1453 -988 -1441 988
rect -1407 -988 -1395 988
rect -1453 -1000 -1395 -988
rect -1275 988 -1217 1000
rect -1275 -988 -1263 988
rect -1229 -988 -1217 988
rect -1275 -1000 -1217 -988
rect -1097 988 -1039 1000
rect -1097 -988 -1085 988
rect -1051 -988 -1039 988
rect -1097 -1000 -1039 -988
rect -919 988 -861 1000
rect -919 -988 -907 988
rect -873 -988 -861 988
rect -919 -1000 -861 -988
rect -741 988 -683 1000
rect -741 -988 -729 988
rect -695 -988 -683 988
rect -741 -1000 -683 -988
rect -563 988 -505 1000
rect -563 -988 -551 988
rect -517 -988 -505 988
rect -563 -1000 -505 -988
rect -385 988 -327 1000
rect -385 -988 -373 988
rect -339 -988 -327 988
rect -385 -1000 -327 -988
rect -207 988 -149 1000
rect -207 -988 -195 988
rect -161 -988 -149 988
rect -207 -1000 -149 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 149 988 207 1000
rect 149 -988 161 988
rect 195 -988 207 988
rect 149 -1000 207 -988
rect 327 988 385 1000
rect 327 -988 339 988
rect 373 -988 385 988
rect 327 -1000 385 -988
rect 505 988 563 1000
rect 505 -988 517 988
rect 551 -988 563 988
rect 505 -1000 563 -988
rect 683 988 741 1000
rect 683 -988 695 988
rect 729 -988 741 988
rect 683 -1000 741 -988
rect 861 988 919 1000
rect 861 -988 873 988
rect 907 -988 919 988
rect 861 -1000 919 -988
rect 1039 988 1097 1000
rect 1039 -988 1051 988
rect 1085 -988 1097 988
rect 1039 -1000 1097 -988
rect 1217 988 1275 1000
rect 1217 -988 1229 988
rect 1263 -988 1275 988
rect 1217 -1000 1275 -988
rect 1395 988 1453 1000
rect 1395 -988 1407 988
rect 1441 -988 1453 988
rect 1395 -1000 1453 -988
rect 1573 988 1631 1000
rect 1573 -988 1585 988
rect 1619 -988 1631 988
rect 1573 -1000 1631 -988
rect 1751 988 1809 1000
rect 1751 -988 1763 988
rect 1797 -988 1809 988
rect 1751 -1000 1809 -988
rect 1929 988 1987 1000
rect 1929 -988 1941 988
rect 1975 -988 1987 988
rect 1929 -1000 1987 -988
rect 2107 988 2165 1000
rect 2107 -988 2119 988
rect 2153 -988 2165 988
rect 2107 -1000 2165 -988
rect 2285 988 2343 1000
rect 2285 -988 2297 988
rect 2331 -988 2343 988
rect 2285 -1000 2343 -988
rect 2463 988 2521 1000
rect 2463 -988 2475 988
rect 2509 -988 2521 988
rect 2463 -1000 2521 -988
rect 2641 988 2699 1000
rect 2641 -988 2653 988
rect 2687 -988 2699 988
rect 2641 -1000 2699 -988
rect 2819 988 2877 1000
rect 2819 -988 2831 988
rect 2865 -988 2877 988
rect 2819 -1000 2877 -988
rect 2997 988 3055 1000
rect 2997 -988 3009 988
rect 3043 -988 3055 988
rect 2997 -1000 3055 -988
rect 3175 988 3233 1000
rect 3175 -988 3187 988
rect 3221 -988 3233 988
rect 3175 -1000 3233 -988
rect 3353 988 3411 1000
rect 3353 -988 3365 988
rect 3399 -988 3411 988
rect 3353 -1000 3411 -988
rect 3531 988 3589 1000
rect 3531 -988 3543 988
rect 3577 -988 3589 988
rect 3531 -1000 3589 -988
rect 3709 988 3767 1000
rect 3709 -988 3721 988
rect 3755 -988 3767 988
rect 3709 -1000 3767 -988
rect 3887 988 3945 1000
rect 3887 -988 3899 988
rect 3933 -988 3945 988
rect 3887 -1000 3945 -988
rect 4065 988 4123 1000
rect 4065 -988 4077 988
rect 4111 -988 4123 988
rect 4065 -1000 4123 -988
rect 4243 988 4301 1000
rect 4243 -988 4255 988
rect 4289 -988 4301 988
rect 4243 -1000 4301 -988
rect 4421 988 4479 1000
rect 4421 -988 4433 988
rect 4467 -988 4479 988
rect 4421 -1000 4479 -988
rect 4599 988 4657 1000
rect 4599 -988 4611 988
rect 4645 -988 4657 988
rect 4599 -1000 4657 -988
rect 4777 988 4835 1000
rect 4777 -988 4789 988
rect 4823 -988 4835 988
rect 4777 -1000 4835 -988
rect 4955 988 5013 1000
rect 4955 -988 4967 988
rect 5001 -988 5013 988
rect 4955 -1000 5013 -988
rect 5133 988 5191 1000
rect 5133 -988 5145 988
rect 5179 -988 5191 988
rect 5133 -1000 5191 -988
rect 5311 988 5369 1000
rect 5311 -988 5323 988
rect 5357 -988 5369 988
rect 5311 -1000 5369 -988
rect 5489 988 5547 1000
rect 5489 -988 5501 988
rect 5535 -988 5547 988
rect 5489 -1000 5547 -988
<< ndiffc >>
rect -5535 -988 -5501 988
rect -5357 -988 -5323 988
rect -5179 -988 -5145 988
rect -5001 -988 -4967 988
rect -4823 -988 -4789 988
rect -4645 -988 -4611 988
rect -4467 -988 -4433 988
rect -4289 -988 -4255 988
rect -4111 -988 -4077 988
rect -3933 -988 -3899 988
rect -3755 -988 -3721 988
rect -3577 -988 -3543 988
rect -3399 -988 -3365 988
rect -3221 -988 -3187 988
rect -3043 -988 -3009 988
rect -2865 -988 -2831 988
rect -2687 -988 -2653 988
rect -2509 -988 -2475 988
rect -2331 -988 -2297 988
rect -2153 -988 -2119 988
rect -1975 -988 -1941 988
rect -1797 -988 -1763 988
rect -1619 -988 -1585 988
rect -1441 -988 -1407 988
rect -1263 -988 -1229 988
rect -1085 -988 -1051 988
rect -907 -988 -873 988
rect -729 -988 -695 988
rect -551 -988 -517 988
rect -373 -988 -339 988
rect -195 -988 -161 988
rect -17 -988 17 988
rect 161 -988 195 988
rect 339 -988 373 988
rect 517 -988 551 988
rect 695 -988 729 988
rect 873 -988 907 988
rect 1051 -988 1085 988
rect 1229 -988 1263 988
rect 1407 -988 1441 988
rect 1585 -988 1619 988
rect 1763 -988 1797 988
rect 1941 -988 1975 988
rect 2119 -988 2153 988
rect 2297 -988 2331 988
rect 2475 -988 2509 988
rect 2653 -988 2687 988
rect 2831 -988 2865 988
rect 3009 -988 3043 988
rect 3187 -988 3221 988
rect 3365 -988 3399 988
rect 3543 -988 3577 988
rect 3721 -988 3755 988
rect 3899 -988 3933 988
rect 4077 -988 4111 988
rect 4255 -988 4289 988
rect 4433 -988 4467 988
rect 4611 -988 4645 988
rect 4789 -988 4823 988
rect 4967 -988 5001 988
rect 5145 -988 5179 988
rect 5323 -988 5357 988
rect 5501 -988 5535 988
<< psubdiff >>
rect -5649 1140 -5553 1174
rect 5553 1140 5649 1174
rect -5649 1078 -5615 1140
rect 5615 1078 5649 1140
rect -5649 -1140 -5615 -1078
rect 5615 -1140 5649 -1078
rect -5649 -1174 -5553 -1140
rect 5553 -1174 5649 -1140
<< psubdiffcont >>
rect -5553 1140 5553 1174
rect -5649 -1078 -5615 1078
rect 5615 -1078 5649 1078
rect -5553 -1174 5553 -1140
<< poly >>
rect -5489 1072 -5369 1088
rect -5489 1038 -5473 1072
rect -5385 1038 -5369 1072
rect -5489 1000 -5369 1038
rect -5311 1072 -5191 1088
rect -5311 1038 -5295 1072
rect -5207 1038 -5191 1072
rect -5311 1000 -5191 1038
rect -5133 1072 -5013 1088
rect -5133 1038 -5117 1072
rect -5029 1038 -5013 1072
rect -5133 1000 -5013 1038
rect -4955 1072 -4835 1088
rect -4955 1038 -4939 1072
rect -4851 1038 -4835 1072
rect -4955 1000 -4835 1038
rect -4777 1072 -4657 1088
rect -4777 1038 -4761 1072
rect -4673 1038 -4657 1072
rect -4777 1000 -4657 1038
rect -4599 1072 -4479 1088
rect -4599 1038 -4583 1072
rect -4495 1038 -4479 1072
rect -4599 1000 -4479 1038
rect -4421 1072 -4301 1088
rect -4421 1038 -4405 1072
rect -4317 1038 -4301 1072
rect -4421 1000 -4301 1038
rect -4243 1072 -4123 1088
rect -4243 1038 -4227 1072
rect -4139 1038 -4123 1072
rect -4243 1000 -4123 1038
rect -4065 1072 -3945 1088
rect -4065 1038 -4049 1072
rect -3961 1038 -3945 1072
rect -4065 1000 -3945 1038
rect -3887 1072 -3767 1088
rect -3887 1038 -3871 1072
rect -3783 1038 -3767 1072
rect -3887 1000 -3767 1038
rect -3709 1072 -3589 1088
rect -3709 1038 -3693 1072
rect -3605 1038 -3589 1072
rect -3709 1000 -3589 1038
rect -3531 1072 -3411 1088
rect -3531 1038 -3515 1072
rect -3427 1038 -3411 1072
rect -3531 1000 -3411 1038
rect -3353 1072 -3233 1088
rect -3353 1038 -3337 1072
rect -3249 1038 -3233 1072
rect -3353 1000 -3233 1038
rect -3175 1072 -3055 1088
rect -3175 1038 -3159 1072
rect -3071 1038 -3055 1072
rect -3175 1000 -3055 1038
rect -2997 1072 -2877 1088
rect -2997 1038 -2981 1072
rect -2893 1038 -2877 1072
rect -2997 1000 -2877 1038
rect -2819 1072 -2699 1088
rect -2819 1038 -2803 1072
rect -2715 1038 -2699 1072
rect -2819 1000 -2699 1038
rect -2641 1072 -2521 1088
rect -2641 1038 -2625 1072
rect -2537 1038 -2521 1072
rect -2641 1000 -2521 1038
rect -2463 1072 -2343 1088
rect -2463 1038 -2447 1072
rect -2359 1038 -2343 1072
rect -2463 1000 -2343 1038
rect -2285 1072 -2165 1088
rect -2285 1038 -2269 1072
rect -2181 1038 -2165 1072
rect -2285 1000 -2165 1038
rect -2107 1072 -1987 1088
rect -2107 1038 -2091 1072
rect -2003 1038 -1987 1072
rect -2107 1000 -1987 1038
rect -1929 1072 -1809 1088
rect -1929 1038 -1913 1072
rect -1825 1038 -1809 1072
rect -1929 1000 -1809 1038
rect -1751 1072 -1631 1088
rect -1751 1038 -1735 1072
rect -1647 1038 -1631 1072
rect -1751 1000 -1631 1038
rect -1573 1072 -1453 1088
rect -1573 1038 -1557 1072
rect -1469 1038 -1453 1072
rect -1573 1000 -1453 1038
rect -1395 1072 -1275 1088
rect -1395 1038 -1379 1072
rect -1291 1038 -1275 1072
rect -1395 1000 -1275 1038
rect -1217 1072 -1097 1088
rect -1217 1038 -1201 1072
rect -1113 1038 -1097 1072
rect -1217 1000 -1097 1038
rect -1039 1072 -919 1088
rect -1039 1038 -1023 1072
rect -935 1038 -919 1072
rect -1039 1000 -919 1038
rect -861 1072 -741 1088
rect -861 1038 -845 1072
rect -757 1038 -741 1072
rect -861 1000 -741 1038
rect -683 1072 -563 1088
rect -683 1038 -667 1072
rect -579 1038 -563 1072
rect -683 1000 -563 1038
rect -505 1072 -385 1088
rect -505 1038 -489 1072
rect -401 1038 -385 1072
rect -505 1000 -385 1038
rect -327 1072 -207 1088
rect -327 1038 -311 1072
rect -223 1038 -207 1072
rect -327 1000 -207 1038
rect -149 1072 -29 1088
rect -149 1038 -133 1072
rect -45 1038 -29 1072
rect -149 1000 -29 1038
rect 29 1072 149 1088
rect 29 1038 45 1072
rect 133 1038 149 1072
rect 29 1000 149 1038
rect 207 1072 327 1088
rect 207 1038 223 1072
rect 311 1038 327 1072
rect 207 1000 327 1038
rect 385 1072 505 1088
rect 385 1038 401 1072
rect 489 1038 505 1072
rect 385 1000 505 1038
rect 563 1072 683 1088
rect 563 1038 579 1072
rect 667 1038 683 1072
rect 563 1000 683 1038
rect 741 1072 861 1088
rect 741 1038 757 1072
rect 845 1038 861 1072
rect 741 1000 861 1038
rect 919 1072 1039 1088
rect 919 1038 935 1072
rect 1023 1038 1039 1072
rect 919 1000 1039 1038
rect 1097 1072 1217 1088
rect 1097 1038 1113 1072
rect 1201 1038 1217 1072
rect 1097 1000 1217 1038
rect 1275 1072 1395 1088
rect 1275 1038 1291 1072
rect 1379 1038 1395 1072
rect 1275 1000 1395 1038
rect 1453 1072 1573 1088
rect 1453 1038 1469 1072
rect 1557 1038 1573 1072
rect 1453 1000 1573 1038
rect 1631 1072 1751 1088
rect 1631 1038 1647 1072
rect 1735 1038 1751 1072
rect 1631 1000 1751 1038
rect 1809 1072 1929 1088
rect 1809 1038 1825 1072
rect 1913 1038 1929 1072
rect 1809 1000 1929 1038
rect 1987 1072 2107 1088
rect 1987 1038 2003 1072
rect 2091 1038 2107 1072
rect 1987 1000 2107 1038
rect 2165 1072 2285 1088
rect 2165 1038 2181 1072
rect 2269 1038 2285 1072
rect 2165 1000 2285 1038
rect 2343 1072 2463 1088
rect 2343 1038 2359 1072
rect 2447 1038 2463 1072
rect 2343 1000 2463 1038
rect 2521 1072 2641 1088
rect 2521 1038 2537 1072
rect 2625 1038 2641 1072
rect 2521 1000 2641 1038
rect 2699 1072 2819 1088
rect 2699 1038 2715 1072
rect 2803 1038 2819 1072
rect 2699 1000 2819 1038
rect 2877 1072 2997 1088
rect 2877 1038 2893 1072
rect 2981 1038 2997 1072
rect 2877 1000 2997 1038
rect 3055 1072 3175 1088
rect 3055 1038 3071 1072
rect 3159 1038 3175 1072
rect 3055 1000 3175 1038
rect 3233 1072 3353 1088
rect 3233 1038 3249 1072
rect 3337 1038 3353 1072
rect 3233 1000 3353 1038
rect 3411 1072 3531 1088
rect 3411 1038 3427 1072
rect 3515 1038 3531 1072
rect 3411 1000 3531 1038
rect 3589 1072 3709 1088
rect 3589 1038 3605 1072
rect 3693 1038 3709 1072
rect 3589 1000 3709 1038
rect 3767 1072 3887 1088
rect 3767 1038 3783 1072
rect 3871 1038 3887 1072
rect 3767 1000 3887 1038
rect 3945 1072 4065 1088
rect 3945 1038 3961 1072
rect 4049 1038 4065 1072
rect 3945 1000 4065 1038
rect 4123 1072 4243 1088
rect 4123 1038 4139 1072
rect 4227 1038 4243 1072
rect 4123 1000 4243 1038
rect 4301 1072 4421 1088
rect 4301 1038 4317 1072
rect 4405 1038 4421 1072
rect 4301 1000 4421 1038
rect 4479 1072 4599 1088
rect 4479 1038 4495 1072
rect 4583 1038 4599 1072
rect 4479 1000 4599 1038
rect 4657 1072 4777 1088
rect 4657 1038 4673 1072
rect 4761 1038 4777 1072
rect 4657 1000 4777 1038
rect 4835 1072 4955 1088
rect 4835 1038 4851 1072
rect 4939 1038 4955 1072
rect 4835 1000 4955 1038
rect 5013 1072 5133 1088
rect 5013 1038 5029 1072
rect 5117 1038 5133 1072
rect 5013 1000 5133 1038
rect 5191 1072 5311 1088
rect 5191 1038 5207 1072
rect 5295 1038 5311 1072
rect 5191 1000 5311 1038
rect 5369 1072 5489 1088
rect 5369 1038 5385 1072
rect 5473 1038 5489 1072
rect 5369 1000 5489 1038
rect -5489 -1038 -5369 -1000
rect -5489 -1072 -5473 -1038
rect -5385 -1072 -5369 -1038
rect -5489 -1088 -5369 -1072
rect -5311 -1038 -5191 -1000
rect -5311 -1072 -5295 -1038
rect -5207 -1072 -5191 -1038
rect -5311 -1088 -5191 -1072
rect -5133 -1038 -5013 -1000
rect -5133 -1072 -5117 -1038
rect -5029 -1072 -5013 -1038
rect -5133 -1088 -5013 -1072
rect -4955 -1038 -4835 -1000
rect -4955 -1072 -4939 -1038
rect -4851 -1072 -4835 -1038
rect -4955 -1088 -4835 -1072
rect -4777 -1038 -4657 -1000
rect -4777 -1072 -4761 -1038
rect -4673 -1072 -4657 -1038
rect -4777 -1088 -4657 -1072
rect -4599 -1038 -4479 -1000
rect -4599 -1072 -4583 -1038
rect -4495 -1072 -4479 -1038
rect -4599 -1088 -4479 -1072
rect -4421 -1038 -4301 -1000
rect -4421 -1072 -4405 -1038
rect -4317 -1072 -4301 -1038
rect -4421 -1088 -4301 -1072
rect -4243 -1038 -4123 -1000
rect -4243 -1072 -4227 -1038
rect -4139 -1072 -4123 -1038
rect -4243 -1088 -4123 -1072
rect -4065 -1038 -3945 -1000
rect -4065 -1072 -4049 -1038
rect -3961 -1072 -3945 -1038
rect -4065 -1088 -3945 -1072
rect -3887 -1038 -3767 -1000
rect -3887 -1072 -3871 -1038
rect -3783 -1072 -3767 -1038
rect -3887 -1088 -3767 -1072
rect -3709 -1038 -3589 -1000
rect -3709 -1072 -3693 -1038
rect -3605 -1072 -3589 -1038
rect -3709 -1088 -3589 -1072
rect -3531 -1038 -3411 -1000
rect -3531 -1072 -3515 -1038
rect -3427 -1072 -3411 -1038
rect -3531 -1088 -3411 -1072
rect -3353 -1038 -3233 -1000
rect -3353 -1072 -3337 -1038
rect -3249 -1072 -3233 -1038
rect -3353 -1088 -3233 -1072
rect -3175 -1038 -3055 -1000
rect -3175 -1072 -3159 -1038
rect -3071 -1072 -3055 -1038
rect -3175 -1088 -3055 -1072
rect -2997 -1038 -2877 -1000
rect -2997 -1072 -2981 -1038
rect -2893 -1072 -2877 -1038
rect -2997 -1088 -2877 -1072
rect -2819 -1038 -2699 -1000
rect -2819 -1072 -2803 -1038
rect -2715 -1072 -2699 -1038
rect -2819 -1088 -2699 -1072
rect -2641 -1038 -2521 -1000
rect -2641 -1072 -2625 -1038
rect -2537 -1072 -2521 -1038
rect -2641 -1088 -2521 -1072
rect -2463 -1038 -2343 -1000
rect -2463 -1072 -2447 -1038
rect -2359 -1072 -2343 -1038
rect -2463 -1088 -2343 -1072
rect -2285 -1038 -2165 -1000
rect -2285 -1072 -2269 -1038
rect -2181 -1072 -2165 -1038
rect -2285 -1088 -2165 -1072
rect -2107 -1038 -1987 -1000
rect -2107 -1072 -2091 -1038
rect -2003 -1072 -1987 -1038
rect -2107 -1088 -1987 -1072
rect -1929 -1038 -1809 -1000
rect -1929 -1072 -1913 -1038
rect -1825 -1072 -1809 -1038
rect -1929 -1088 -1809 -1072
rect -1751 -1038 -1631 -1000
rect -1751 -1072 -1735 -1038
rect -1647 -1072 -1631 -1038
rect -1751 -1088 -1631 -1072
rect -1573 -1038 -1453 -1000
rect -1573 -1072 -1557 -1038
rect -1469 -1072 -1453 -1038
rect -1573 -1088 -1453 -1072
rect -1395 -1038 -1275 -1000
rect -1395 -1072 -1379 -1038
rect -1291 -1072 -1275 -1038
rect -1395 -1088 -1275 -1072
rect -1217 -1038 -1097 -1000
rect -1217 -1072 -1201 -1038
rect -1113 -1072 -1097 -1038
rect -1217 -1088 -1097 -1072
rect -1039 -1038 -919 -1000
rect -1039 -1072 -1023 -1038
rect -935 -1072 -919 -1038
rect -1039 -1088 -919 -1072
rect -861 -1038 -741 -1000
rect -861 -1072 -845 -1038
rect -757 -1072 -741 -1038
rect -861 -1088 -741 -1072
rect -683 -1038 -563 -1000
rect -683 -1072 -667 -1038
rect -579 -1072 -563 -1038
rect -683 -1088 -563 -1072
rect -505 -1038 -385 -1000
rect -505 -1072 -489 -1038
rect -401 -1072 -385 -1038
rect -505 -1088 -385 -1072
rect -327 -1038 -207 -1000
rect -327 -1072 -311 -1038
rect -223 -1072 -207 -1038
rect -327 -1088 -207 -1072
rect -149 -1038 -29 -1000
rect -149 -1072 -133 -1038
rect -45 -1072 -29 -1038
rect -149 -1088 -29 -1072
rect 29 -1038 149 -1000
rect 29 -1072 45 -1038
rect 133 -1072 149 -1038
rect 29 -1088 149 -1072
rect 207 -1038 327 -1000
rect 207 -1072 223 -1038
rect 311 -1072 327 -1038
rect 207 -1088 327 -1072
rect 385 -1038 505 -1000
rect 385 -1072 401 -1038
rect 489 -1072 505 -1038
rect 385 -1088 505 -1072
rect 563 -1038 683 -1000
rect 563 -1072 579 -1038
rect 667 -1072 683 -1038
rect 563 -1088 683 -1072
rect 741 -1038 861 -1000
rect 741 -1072 757 -1038
rect 845 -1072 861 -1038
rect 741 -1088 861 -1072
rect 919 -1038 1039 -1000
rect 919 -1072 935 -1038
rect 1023 -1072 1039 -1038
rect 919 -1088 1039 -1072
rect 1097 -1038 1217 -1000
rect 1097 -1072 1113 -1038
rect 1201 -1072 1217 -1038
rect 1097 -1088 1217 -1072
rect 1275 -1038 1395 -1000
rect 1275 -1072 1291 -1038
rect 1379 -1072 1395 -1038
rect 1275 -1088 1395 -1072
rect 1453 -1038 1573 -1000
rect 1453 -1072 1469 -1038
rect 1557 -1072 1573 -1038
rect 1453 -1088 1573 -1072
rect 1631 -1038 1751 -1000
rect 1631 -1072 1647 -1038
rect 1735 -1072 1751 -1038
rect 1631 -1088 1751 -1072
rect 1809 -1038 1929 -1000
rect 1809 -1072 1825 -1038
rect 1913 -1072 1929 -1038
rect 1809 -1088 1929 -1072
rect 1987 -1038 2107 -1000
rect 1987 -1072 2003 -1038
rect 2091 -1072 2107 -1038
rect 1987 -1088 2107 -1072
rect 2165 -1038 2285 -1000
rect 2165 -1072 2181 -1038
rect 2269 -1072 2285 -1038
rect 2165 -1088 2285 -1072
rect 2343 -1038 2463 -1000
rect 2343 -1072 2359 -1038
rect 2447 -1072 2463 -1038
rect 2343 -1088 2463 -1072
rect 2521 -1038 2641 -1000
rect 2521 -1072 2537 -1038
rect 2625 -1072 2641 -1038
rect 2521 -1088 2641 -1072
rect 2699 -1038 2819 -1000
rect 2699 -1072 2715 -1038
rect 2803 -1072 2819 -1038
rect 2699 -1088 2819 -1072
rect 2877 -1038 2997 -1000
rect 2877 -1072 2893 -1038
rect 2981 -1072 2997 -1038
rect 2877 -1088 2997 -1072
rect 3055 -1038 3175 -1000
rect 3055 -1072 3071 -1038
rect 3159 -1072 3175 -1038
rect 3055 -1088 3175 -1072
rect 3233 -1038 3353 -1000
rect 3233 -1072 3249 -1038
rect 3337 -1072 3353 -1038
rect 3233 -1088 3353 -1072
rect 3411 -1038 3531 -1000
rect 3411 -1072 3427 -1038
rect 3515 -1072 3531 -1038
rect 3411 -1088 3531 -1072
rect 3589 -1038 3709 -1000
rect 3589 -1072 3605 -1038
rect 3693 -1072 3709 -1038
rect 3589 -1088 3709 -1072
rect 3767 -1038 3887 -1000
rect 3767 -1072 3783 -1038
rect 3871 -1072 3887 -1038
rect 3767 -1088 3887 -1072
rect 3945 -1038 4065 -1000
rect 3945 -1072 3961 -1038
rect 4049 -1072 4065 -1038
rect 3945 -1088 4065 -1072
rect 4123 -1038 4243 -1000
rect 4123 -1072 4139 -1038
rect 4227 -1072 4243 -1038
rect 4123 -1088 4243 -1072
rect 4301 -1038 4421 -1000
rect 4301 -1072 4317 -1038
rect 4405 -1072 4421 -1038
rect 4301 -1088 4421 -1072
rect 4479 -1038 4599 -1000
rect 4479 -1072 4495 -1038
rect 4583 -1072 4599 -1038
rect 4479 -1088 4599 -1072
rect 4657 -1038 4777 -1000
rect 4657 -1072 4673 -1038
rect 4761 -1072 4777 -1038
rect 4657 -1088 4777 -1072
rect 4835 -1038 4955 -1000
rect 4835 -1072 4851 -1038
rect 4939 -1072 4955 -1038
rect 4835 -1088 4955 -1072
rect 5013 -1038 5133 -1000
rect 5013 -1072 5029 -1038
rect 5117 -1072 5133 -1038
rect 5013 -1088 5133 -1072
rect 5191 -1038 5311 -1000
rect 5191 -1072 5207 -1038
rect 5295 -1072 5311 -1038
rect 5191 -1088 5311 -1072
rect 5369 -1038 5489 -1000
rect 5369 -1072 5385 -1038
rect 5473 -1072 5489 -1038
rect 5369 -1088 5489 -1072
<< polycont >>
rect -5473 1038 -5385 1072
rect -5295 1038 -5207 1072
rect -5117 1038 -5029 1072
rect -4939 1038 -4851 1072
rect -4761 1038 -4673 1072
rect -4583 1038 -4495 1072
rect -4405 1038 -4317 1072
rect -4227 1038 -4139 1072
rect -4049 1038 -3961 1072
rect -3871 1038 -3783 1072
rect -3693 1038 -3605 1072
rect -3515 1038 -3427 1072
rect -3337 1038 -3249 1072
rect -3159 1038 -3071 1072
rect -2981 1038 -2893 1072
rect -2803 1038 -2715 1072
rect -2625 1038 -2537 1072
rect -2447 1038 -2359 1072
rect -2269 1038 -2181 1072
rect -2091 1038 -2003 1072
rect -1913 1038 -1825 1072
rect -1735 1038 -1647 1072
rect -1557 1038 -1469 1072
rect -1379 1038 -1291 1072
rect -1201 1038 -1113 1072
rect -1023 1038 -935 1072
rect -845 1038 -757 1072
rect -667 1038 -579 1072
rect -489 1038 -401 1072
rect -311 1038 -223 1072
rect -133 1038 -45 1072
rect 45 1038 133 1072
rect 223 1038 311 1072
rect 401 1038 489 1072
rect 579 1038 667 1072
rect 757 1038 845 1072
rect 935 1038 1023 1072
rect 1113 1038 1201 1072
rect 1291 1038 1379 1072
rect 1469 1038 1557 1072
rect 1647 1038 1735 1072
rect 1825 1038 1913 1072
rect 2003 1038 2091 1072
rect 2181 1038 2269 1072
rect 2359 1038 2447 1072
rect 2537 1038 2625 1072
rect 2715 1038 2803 1072
rect 2893 1038 2981 1072
rect 3071 1038 3159 1072
rect 3249 1038 3337 1072
rect 3427 1038 3515 1072
rect 3605 1038 3693 1072
rect 3783 1038 3871 1072
rect 3961 1038 4049 1072
rect 4139 1038 4227 1072
rect 4317 1038 4405 1072
rect 4495 1038 4583 1072
rect 4673 1038 4761 1072
rect 4851 1038 4939 1072
rect 5029 1038 5117 1072
rect 5207 1038 5295 1072
rect 5385 1038 5473 1072
rect -5473 -1072 -5385 -1038
rect -5295 -1072 -5207 -1038
rect -5117 -1072 -5029 -1038
rect -4939 -1072 -4851 -1038
rect -4761 -1072 -4673 -1038
rect -4583 -1072 -4495 -1038
rect -4405 -1072 -4317 -1038
rect -4227 -1072 -4139 -1038
rect -4049 -1072 -3961 -1038
rect -3871 -1072 -3783 -1038
rect -3693 -1072 -3605 -1038
rect -3515 -1072 -3427 -1038
rect -3337 -1072 -3249 -1038
rect -3159 -1072 -3071 -1038
rect -2981 -1072 -2893 -1038
rect -2803 -1072 -2715 -1038
rect -2625 -1072 -2537 -1038
rect -2447 -1072 -2359 -1038
rect -2269 -1072 -2181 -1038
rect -2091 -1072 -2003 -1038
rect -1913 -1072 -1825 -1038
rect -1735 -1072 -1647 -1038
rect -1557 -1072 -1469 -1038
rect -1379 -1072 -1291 -1038
rect -1201 -1072 -1113 -1038
rect -1023 -1072 -935 -1038
rect -845 -1072 -757 -1038
rect -667 -1072 -579 -1038
rect -489 -1072 -401 -1038
rect -311 -1072 -223 -1038
rect -133 -1072 -45 -1038
rect 45 -1072 133 -1038
rect 223 -1072 311 -1038
rect 401 -1072 489 -1038
rect 579 -1072 667 -1038
rect 757 -1072 845 -1038
rect 935 -1072 1023 -1038
rect 1113 -1072 1201 -1038
rect 1291 -1072 1379 -1038
rect 1469 -1072 1557 -1038
rect 1647 -1072 1735 -1038
rect 1825 -1072 1913 -1038
rect 2003 -1072 2091 -1038
rect 2181 -1072 2269 -1038
rect 2359 -1072 2447 -1038
rect 2537 -1072 2625 -1038
rect 2715 -1072 2803 -1038
rect 2893 -1072 2981 -1038
rect 3071 -1072 3159 -1038
rect 3249 -1072 3337 -1038
rect 3427 -1072 3515 -1038
rect 3605 -1072 3693 -1038
rect 3783 -1072 3871 -1038
rect 3961 -1072 4049 -1038
rect 4139 -1072 4227 -1038
rect 4317 -1072 4405 -1038
rect 4495 -1072 4583 -1038
rect 4673 -1072 4761 -1038
rect 4851 -1072 4939 -1038
rect 5029 -1072 5117 -1038
rect 5207 -1072 5295 -1038
rect 5385 -1072 5473 -1038
<< locali >>
rect -5649 1140 -5553 1174
rect 5553 1140 5649 1174
rect -5649 1078 -5615 1140
rect 5615 1078 5649 1140
rect -5489 1038 -5473 1072
rect -5385 1038 -5369 1072
rect -5311 1038 -5295 1072
rect -5207 1038 -5191 1072
rect -5133 1038 -5117 1072
rect -5029 1038 -5013 1072
rect -4955 1038 -4939 1072
rect -4851 1038 -4835 1072
rect -4777 1038 -4761 1072
rect -4673 1038 -4657 1072
rect -4599 1038 -4583 1072
rect -4495 1038 -4479 1072
rect -4421 1038 -4405 1072
rect -4317 1038 -4301 1072
rect -4243 1038 -4227 1072
rect -4139 1038 -4123 1072
rect -4065 1038 -4049 1072
rect -3961 1038 -3945 1072
rect -3887 1038 -3871 1072
rect -3783 1038 -3767 1072
rect -3709 1038 -3693 1072
rect -3605 1038 -3589 1072
rect -3531 1038 -3515 1072
rect -3427 1038 -3411 1072
rect -3353 1038 -3337 1072
rect -3249 1038 -3233 1072
rect -3175 1038 -3159 1072
rect -3071 1038 -3055 1072
rect -2997 1038 -2981 1072
rect -2893 1038 -2877 1072
rect -2819 1038 -2803 1072
rect -2715 1038 -2699 1072
rect -2641 1038 -2625 1072
rect -2537 1038 -2521 1072
rect -2463 1038 -2447 1072
rect -2359 1038 -2343 1072
rect -2285 1038 -2269 1072
rect -2181 1038 -2165 1072
rect -2107 1038 -2091 1072
rect -2003 1038 -1987 1072
rect -1929 1038 -1913 1072
rect -1825 1038 -1809 1072
rect -1751 1038 -1735 1072
rect -1647 1038 -1631 1072
rect -1573 1038 -1557 1072
rect -1469 1038 -1453 1072
rect -1395 1038 -1379 1072
rect -1291 1038 -1275 1072
rect -1217 1038 -1201 1072
rect -1113 1038 -1097 1072
rect -1039 1038 -1023 1072
rect -935 1038 -919 1072
rect -861 1038 -845 1072
rect -757 1038 -741 1072
rect -683 1038 -667 1072
rect -579 1038 -563 1072
rect -505 1038 -489 1072
rect -401 1038 -385 1072
rect -327 1038 -311 1072
rect -223 1038 -207 1072
rect -149 1038 -133 1072
rect -45 1038 -29 1072
rect 29 1038 45 1072
rect 133 1038 149 1072
rect 207 1038 223 1072
rect 311 1038 327 1072
rect 385 1038 401 1072
rect 489 1038 505 1072
rect 563 1038 579 1072
rect 667 1038 683 1072
rect 741 1038 757 1072
rect 845 1038 861 1072
rect 919 1038 935 1072
rect 1023 1038 1039 1072
rect 1097 1038 1113 1072
rect 1201 1038 1217 1072
rect 1275 1038 1291 1072
rect 1379 1038 1395 1072
rect 1453 1038 1469 1072
rect 1557 1038 1573 1072
rect 1631 1038 1647 1072
rect 1735 1038 1751 1072
rect 1809 1038 1825 1072
rect 1913 1038 1929 1072
rect 1987 1038 2003 1072
rect 2091 1038 2107 1072
rect 2165 1038 2181 1072
rect 2269 1038 2285 1072
rect 2343 1038 2359 1072
rect 2447 1038 2463 1072
rect 2521 1038 2537 1072
rect 2625 1038 2641 1072
rect 2699 1038 2715 1072
rect 2803 1038 2819 1072
rect 2877 1038 2893 1072
rect 2981 1038 2997 1072
rect 3055 1038 3071 1072
rect 3159 1038 3175 1072
rect 3233 1038 3249 1072
rect 3337 1038 3353 1072
rect 3411 1038 3427 1072
rect 3515 1038 3531 1072
rect 3589 1038 3605 1072
rect 3693 1038 3709 1072
rect 3767 1038 3783 1072
rect 3871 1038 3887 1072
rect 3945 1038 3961 1072
rect 4049 1038 4065 1072
rect 4123 1038 4139 1072
rect 4227 1038 4243 1072
rect 4301 1038 4317 1072
rect 4405 1038 4421 1072
rect 4479 1038 4495 1072
rect 4583 1038 4599 1072
rect 4657 1038 4673 1072
rect 4761 1038 4777 1072
rect 4835 1038 4851 1072
rect 4939 1038 4955 1072
rect 5013 1038 5029 1072
rect 5117 1038 5133 1072
rect 5191 1038 5207 1072
rect 5295 1038 5311 1072
rect 5369 1038 5385 1072
rect 5473 1038 5489 1072
rect -5535 988 -5501 1004
rect -5535 -1004 -5501 -988
rect -5357 988 -5323 1004
rect -5357 -1004 -5323 -988
rect -5179 988 -5145 1004
rect -5179 -1004 -5145 -988
rect -5001 988 -4967 1004
rect -5001 -1004 -4967 -988
rect -4823 988 -4789 1004
rect -4823 -1004 -4789 -988
rect -4645 988 -4611 1004
rect -4645 -1004 -4611 -988
rect -4467 988 -4433 1004
rect -4467 -1004 -4433 -988
rect -4289 988 -4255 1004
rect -4289 -1004 -4255 -988
rect -4111 988 -4077 1004
rect -4111 -1004 -4077 -988
rect -3933 988 -3899 1004
rect -3933 -1004 -3899 -988
rect -3755 988 -3721 1004
rect -3755 -1004 -3721 -988
rect -3577 988 -3543 1004
rect -3577 -1004 -3543 -988
rect -3399 988 -3365 1004
rect -3399 -1004 -3365 -988
rect -3221 988 -3187 1004
rect -3221 -1004 -3187 -988
rect -3043 988 -3009 1004
rect -3043 -1004 -3009 -988
rect -2865 988 -2831 1004
rect -2865 -1004 -2831 -988
rect -2687 988 -2653 1004
rect -2687 -1004 -2653 -988
rect -2509 988 -2475 1004
rect -2509 -1004 -2475 -988
rect -2331 988 -2297 1004
rect -2331 -1004 -2297 -988
rect -2153 988 -2119 1004
rect -2153 -1004 -2119 -988
rect -1975 988 -1941 1004
rect -1975 -1004 -1941 -988
rect -1797 988 -1763 1004
rect -1797 -1004 -1763 -988
rect -1619 988 -1585 1004
rect -1619 -1004 -1585 -988
rect -1441 988 -1407 1004
rect -1441 -1004 -1407 -988
rect -1263 988 -1229 1004
rect -1263 -1004 -1229 -988
rect -1085 988 -1051 1004
rect -1085 -1004 -1051 -988
rect -907 988 -873 1004
rect -907 -1004 -873 -988
rect -729 988 -695 1004
rect -729 -1004 -695 -988
rect -551 988 -517 1004
rect -551 -1004 -517 -988
rect -373 988 -339 1004
rect -373 -1004 -339 -988
rect -195 988 -161 1004
rect -195 -1004 -161 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 161 988 195 1004
rect 161 -1004 195 -988
rect 339 988 373 1004
rect 339 -1004 373 -988
rect 517 988 551 1004
rect 517 -1004 551 -988
rect 695 988 729 1004
rect 695 -1004 729 -988
rect 873 988 907 1004
rect 873 -1004 907 -988
rect 1051 988 1085 1004
rect 1051 -1004 1085 -988
rect 1229 988 1263 1004
rect 1229 -1004 1263 -988
rect 1407 988 1441 1004
rect 1407 -1004 1441 -988
rect 1585 988 1619 1004
rect 1585 -1004 1619 -988
rect 1763 988 1797 1004
rect 1763 -1004 1797 -988
rect 1941 988 1975 1004
rect 1941 -1004 1975 -988
rect 2119 988 2153 1004
rect 2119 -1004 2153 -988
rect 2297 988 2331 1004
rect 2297 -1004 2331 -988
rect 2475 988 2509 1004
rect 2475 -1004 2509 -988
rect 2653 988 2687 1004
rect 2653 -1004 2687 -988
rect 2831 988 2865 1004
rect 2831 -1004 2865 -988
rect 3009 988 3043 1004
rect 3009 -1004 3043 -988
rect 3187 988 3221 1004
rect 3187 -1004 3221 -988
rect 3365 988 3399 1004
rect 3365 -1004 3399 -988
rect 3543 988 3577 1004
rect 3543 -1004 3577 -988
rect 3721 988 3755 1004
rect 3721 -1004 3755 -988
rect 3899 988 3933 1004
rect 3899 -1004 3933 -988
rect 4077 988 4111 1004
rect 4077 -1004 4111 -988
rect 4255 988 4289 1004
rect 4255 -1004 4289 -988
rect 4433 988 4467 1004
rect 4433 -1004 4467 -988
rect 4611 988 4645 1004
rect 4611 -1004 4645 -988
rect 4789 988 4823 1004
rect 4789 -1004 4823 -988
rect 4967 988 5001 1004
rect 4967 -1004 5001 -988
rect 5145 988 5179 1004
rect 5145 -1004 5179 -988
rect 5323 988 5357 1004
rect 5323 -1004 5357 -988
rect 5501 988 5535 1004
rect 5501 -1004 5535 -988
rect -5489 -1072 -5473 -1038
rect -5385 -1072 -5369 -1038
rect -5311 -1072 -5295 -1038
rect -5207 -1072 -5191 -1038
rect -5133 -1072 -5117 -1038
rect -5029 -1072 -5013 -1038
rect -4955 -1072 -4939 -1038
rect -4851 -1072 -4835 -1038
rect -4777 -1072 -4761 -1038
rect -4673 -1072 -4657 -1038
rect -4599 -1072 -4583 -1038
rect -4495 -1072 -4479 -1038
rect -4421 -1072 -4405 -1038
rect -4317 -1072 -4301 -1038
rect -4243 -1072 -4227 -1038
rect -4139 -1072 -4123 -1038
rect -4065 -1072 -4049 -1038
rect -3961 -1072 -3945 -1038
rect -3887 -1072 -3871 -1038
rect -3783 -1072 -3767 -1038
rect -3709 -1072 -3693 -1038
rect -3605 -1072 -3589 -1038
rect -3531 -1072 -3515 -1038
rect -3427 -1072 -3411 -1038
rect -3353 -1072 -3337 -1038
rect -3249 -1072 -3233 -1038
rect -3175 -1072 -3159 -1038
rect -3071 -1072 -3055 -1038
rect -2997 -1072 -2981 -1038
rect -2893 -1072 -2877 -1038
rect -2819 -1072 -2803 -1038
rect -2715 -1072 -2699 -1038
rect -2641 -1072 -2625 -1038
rect -2537 -1072 -2521 -1038
rect -2463 -1072 -2447 -1038
rect -2359 -1072 -2343 -1038
rect -2285 -1072 -2269 -1038
rect -2181 -1072 -2165 -1038
rect -2107 -1072 -2091 -1038
rect -2003 -1072 -1987 -1038
rect -1929 -1072 -1913 -1038
rect -1825 -1072 -1809 -1038
rect -1751 -1072 -1735 -1038
rect -1647 -1072 -1631 -1038
rect -1573 -1072 -1557 -1038
rect -1469 -1072 -1453 -1038
rect -1395 -1072 -1379 -1038
rect -1291 -1072 -1275 -1038
rect -1217 -1072 -1201 -1038
rect -1113 -1072 -1097 -1038
rect -1039 -1072 -1023 -1038
rect -935 -1072 -919 -1038
rect -861 -1072 -845 -1038
rect -757 -1072 -741 -1038
rect -683 -1072 -667 -1038
rect -579 -1072 -563 -1038
rect -505 -1072 -489 -1038
rect -401 -1072 -385 -1038
rect -327 -1072 -311 -1038
rect -223 -1072 -207 -1038
rect -149 -1072 -133 -1038
rect -45 -1072 -29 -1038
rect 29 -1072 45 -1038
rect 133 -1072 149 -1038
rect 207 -1072 223 -1038
rect 311 -1072 327 -1038
rect 385 -1072 401 -1038
rect 489 -1072 505 -1038
rect 563 -1072 579 -1038
rect 667 -1072 683 -1038
rect 741 -1072 757 -1038
rect 845 -1072 861 -1038
rect 919 -1072 935 -1038
rect 1023 -1072 1039 -1038
rect 1097 -1072 1113 -1038
rect 1201 -1072 1217 -1038
rect 1275 -1072 1291 -1038
rect 1379 -1072 1395 -1038
rect 1453 -1072 1469 -1038
rect 1557 -1072 1573 -1038
rect 1631 -1072 1647 -1038
rect 1735 -1072 1751 -1038
rect 1809 -1072 1825 -1038
rect 1913 -1072 1929 -1038
rect 1987 -1072 2003 -1038
rect 2091 -1072 2107 -1038
rect 2165 -1072 2181 -1038
rect 2269 -1072 2285 -1038
rect 2343 -1072 2359 -1038
rect 2447 -1072 2463 -1038
rect 2521 -1072 2537 -1038
rect 2625 -1072 2641 -1038
rect 2699 -1072 2715 -1038
rect 2803 -1072 2819 -1038
rect 2877 -1072 2893 -1038
rect 2981 -1072 2997 -1038
rect 3055 -1072 3071 -1038
rect 3159 -1072 3175 -1038
rect 3233 -1072 3249 -1038
rect 3337 -1072 3353 -1038
rect 3411 -1072 3427 -1038
rect 3515 -1072 3531 -1038
rect 3589 -1072 3605 -1038
rect 3693 -1072 3709 -1038
rect 3767 -1072 3783 -1038
rect 3871 -1072 3887 -1038
rect 3945 -1072 3961 -1038
rect 4049 -1072 4065 -1038
rect 4123 -1072 4139 -1038
rect 4227 -1072 4243 -1038
rect 4301 -1072 4317 -1038
rect 4405 -1072 4421 -1038
rect 4479 -1072 4495 -1038
rect 4583 -1072 4599 -1038
rect 4657 -1072 4673 -1038
rect 4761 -1072 4777 -1038
rect 4835 -1072 4851 -1038
rect 4939 -1072 4955 -1038
rect 5013 -1072 5029 -1038
rect 5117 -1072 5133 -1038
rect 5191 -1072 5207 -1038
rect 5295 -1072 5311 -1038
rect 5369 -1072 5385 -1038
rect 5473 -1072 5489 -1038
rect -5649 -1140 -5615 -1078
rect 5615 -1140 5649 -1078
rect -5649 -1174 -5553 -1140
rect 5553 -1174 5649 -1140
<< viali >>
rect -5473 1038 -5385 1072
rect -5295 1038 -5207 1072
rect -5117 1038 -5029 1072
rect -4939 1038 -4851 1072
rect -4761 1038 -4673 1072
rect -4583 1038 -4495 1072
rect -4405 1038 -4317 1072
rect -4227 1038 -4139 1072
rect -4049 1038 -3961 1072
rect -3871 1038 -3783 1072
rect -3693 1038 -3605 1072
rect -3515 1038 -3427 1072
rect -3337 1038 -3249 1072
rect -3159 1038 -3071 1072
rect -2981 1038 -2893 1072
rect -2803 1038 -2715 1072
rect -2625 1038 -2537 1072
rect -2447 1038 -2359 1072
rect -2269 1038 -2181 1072
rect -2091 1038 -2003 1072
rect -1913 1038 -1825 1072
rect -1735 1038 -1647 1072
rect -1557 1038 -1469 1072
rect -1379 1038 -1291 1072
rect -1201 1038 -1113 1072
rect -1023 1038 -935 1072
rect -845 1038 -757 1072
rect -667 1038 -579 1072
rect -489 1038 -401 1072
rect -311 1038 -223 1072
rect -133 1038 -45 1072
rect 45 1038 133 1072
rect 223 1038 311 1072
rect 401 1038 489 1072
rect 579 1038 667 1072
rect 757 1038 845 1072
rect 935 1038 1023 1072
rect 1113 1038 1201 1072
rect 1291 1038 1379 1072
rect 1469 1038 1557 1072
rect 1647 1038 1735 1072
rect 1825 1038 1913 1072
rect 2003 1038 2091 1072
rect 2181 1038 2269 1072
rect 2359 1038 2447 1072
rect 2537 1038 2625 1072
rect 2715 1038 2803 1072
rect 2893 1038 2981 1072
rect 3071 1038 3159 1072
rect 3249 1038 3337 1072
rect 3427 1038 3515 1072
rect 3605 1038 3693 1072
rect 3783 1038 3871 1072
rect 3961 1038 4049 1072
rect 4139 1038 4227 1072
rect 4317 1038 4405 1072
rect 4495 1038 4583 1072
rect 4673 1038 4761 1072
rect 4851 1038 4939 1072
rect 5029 1038 5117 1072
rect 5207 1038 5295 1072
rect 5385 1038 5473 1072
rect -5535 -988 -5501 988
rect -5357 -988 -5323 988
rect -5179 -988 -5145 988
rect -5001 -988 -4967 988
rect -4823 -988 -4789 988
rect -4645 -988 -4611 988
rect -4467 -988 -4433 988
rect -4289 -988 -4255 988
rect -4111 -988 -4077 988
rect -3933 -988 -3899 988
rect -3755 -988 -3721 988
rect -3577 -988 -3543 988
rect -3399 -988 -3365 988
rect -3221 -988 -3187 988
rect -3043 -988 -3009 988
rect -2865 -988 -2831 988
rect -2687 -988 -2653 988
rect -2509 -988 -2475 988
rect -2331 -988 -2297 988
rect -2153 -988 -2119 988
rect -1975 -988 -1941 988
rect -1797 -988 -1763 988
rect -1619 -988 -1585 988
rect -1441 -988 -1407 988
rect -1263 -988 -1229 988
rect -1085 -988 -1051 988
rect -907 -988 -873 988
rect -729 -988 -695 988
rect -551 -988 -517 988
rect -373 -988 -339 988
rect -195 -988 -161 988
rect -17 -988 17 988
rect 161 -988 195 988
rect 339 -988 373 988
rect 517 -988 551 988
rect 695 -988 729 988
rect 873 -988 907 988
rect 1051 -988 1085 988
rect 1229 -988 1263 988
rect 1407 -988 1441 988
rect 1585 -988 1619 988
rect 1763 -988 1797 988
rect 1941 -988 1975 988
rect 2119 -988 2153 988
rect 2297 -988 2331 988
rect 2475 -988 2509 988
rect 2653 -988 2687 988
rect 2831 -988 2865 988
rect 3009 -988 3043 988
rect 3187 -988 3221 988
rect 3365 -988 3399 988
rect 3543 -988 3577 988
rect 3721 -988 3755 988
rect 3899 -988 3933 988
rect 4077 -988 4111 988
rect 4255 -988 4289 988
rect 4433 -988 4467 988
rect 4611 -988 4645 988
rect 4789 -988 4823 988
rect 4967 -988 5001 988
rect 5145 -988 5179 988
rect 5323 -988 5357 988
rect 5501 -988 5535 988
rect -5473 -1072 -5385 -1038
rect -5295 -1072 -5207 -1038
rect -5117 -1072 -5029 -1038
rect -4939 -1072 -4851 -1038
rect -4761 -1072 -4673 -1038
rect -4583 -1072 -4495 -1038
rect -4405 -1072 -4317 -1038
rect -4227 -1072 -4139 -1038
rect -4049 -1072 -3961 -1038
rect -3871 -1072 -3783 -1038
rect -3693 -1072 -3605 -1038
rect -3515 -1072 -3427 -1038
rect -3337 -1072 -3249 -1038
rect -3159 -1072 -3071 -1038
rect -2981 -1072 -2893 -1038
rect -2803 -1072 -2715 -1038
rect -2625 -1072 -2537 -1038
rect -2447 -1072 -2359 -1038
rect -2269 -1072 -2181 -1038
rect -2091 -1072 -2003 -1038
rect -1913 -1072 -1825 -1038
rect -1735 -1072 -1647 -1038
rect -1557 -1072 -1469 -1038
rect -1379 -1072 -1291 -1038
rect -1201 -1072 -1113 -1038
rect -1023 -1072 -935 -1038
rect -845 -1072 -757 -1038
rect -667 -1072 -579 -1038
rect -489 -1072 -401 -1038
rect -311 -1072 -223 -1038
rect -133 -1072 -45 -1038
rect 45 -1072 133 -1038
rect 223 -1072 311 -1038
rect 401 -1072 489 -1038
rect 579 -1072 667 -1038
rect 757 -1072 845 -1038
rect 935 -1072 1023 -1038
rect 1113 -1072 1201 -1038
rect 1291 -1072 1379 -1038
rect 1469 -1072 1557 -1038
rect 1647 -1072 1735 -1038
rect 1825 -1072 1913 -1038
rect 2003 -1072 2091 -1038
rect 2181 -1072 2269 -1038
rect 2359 -1072 2447 -1038
rect 2537 -1072 2625 -1038
rect 2715 -1072 2803 -1038
rect 2893 -1072 2981 -1038
rect 3071 -1072 3159 -1038
rect 3249 -1072 3337 -1038
rect 3427 -1072 3515 -1038
rect 3605 -1072 3693 -1038
rect 3783 -1072 3871 -1038
rect 3961 -1072 4049 -1038
rect 4139 -1072 4227 -1038
rect 4317 -1072 4405 -1038
rect 4495 -1072 4583 -1038
rect 4673 -1072 4761 -1038
rect 4851 -1072 4939 -1038
rect 5029 -1072 5117 -1038
rect 5207 -1072 5295 -1038
rect 5385 -1072 5473 -1038
<< metal1 >>
rect -5485 1072 -5373 1078
rect -5485 1038 -5473 1072
rect -5385 1038 -5373 1072
rect -5485 1032 -5373 1038
rect -5307 1072 -5195 1078
rect -5307 1038 -5295 1072
rect -5207 1038 -5195 1072
rect -5307 1032 -5195 1038
rect -5129 1072 -5017 1078
rect -5129 1038 -5117 1072
rect -5029 1038 -5017 1072
rect -5129 1032 -5017 1038
rect -4951 1072 -4839 1078
rect -4951 1038 -4939 1072
rect -4851 1038 -4839 1072
rect -4951 1032 -4839 1038
rect -4773 1072 -4661 1078
rect -4773 1038 -4761 1072
rect -4673 1038 -4661 1072
rect -4773 1032 -4661 1038
rect -4595 1072 -4483 1078
rect -4595 1038 -4583 1072
rect -4495 1038 -4483 1072
rect -4595 1032 -4483 1038
rect -4417 1072 -4305 1078
rect -4417 1038 -4405 1072
rect -4317 1038 -4305 1072
rect -4417 1032 -4305 1038
rect -4239 1072 -4127 1078
rect -4239 1038 -4227 1072
rect -4139 1038 -4127 1072
rect -4239 1032 -4127 1038
rect -4061 1072 -3949 1078
rect -4061 1038 -4049 1072
rect -3961 1038 -3949 1072
rect -4061 1032 -3949 1038
rect -3883 1072 -3771 1078
rect -3883 1038 -3871 1072
rect -3783 1038 -3771 1072
rect -3883 1032 -3771 1038
rect -3705 1072 -3593 1078
rect -3705 1038 -3693 1072
rect -3605 1038 -3593 1072
rect -3705 1032 -3593 1038
rect -3527 1072 -3415 1078
rect -3527 1038 -3515 1072
rect -3427 1038 -3415 1072
rect -3527 1032 -3415 1038
rect -3349 1072 -3237 1078
rect -3349 1038 -3337 1072
rect -3249 1038 -3237 1072
rect -3349 1032 -3237 1038
rect -3171 1072 -3059 1078
rect -3171 1038 -3159 1072
rect -3071 1038 -3059 1072
rect -3171 1032 -3059 1038
rect -2993 1072 -2881 1078
rect -2993 1038 -2981 1072
rect -2893 1038 -2881 1072
rect -2993 1032 -2881 1038
rect -2815 1072 -2703 1078
rect -2815 1038 -2803 1072
rect -2715 1038 -2703 1072
rect -2815 1032 -2703 1038
rect -2637 1072 -2525 1078
rect -2637 1038 -2625 1072
rect -2537 1038 -2525 1072
rect -2637 1032 -2525 1038
rect -2459 1072 -2347 1078
rect -2459 1038 -2447 1072
rect -2359 1038 -2347 1072
rect -2459 1032 -2347 1038
rect -2281 1072 -2169 1078
rect -2281 1038 -2269 1072
rect -2181 1038 -2169 1072
rect -2281 1032 -2169 1038
rect -2103 1072 -1991 1078
rect -2103 1038 -2091 1072
rect -2003 1038 -1991 1072
rect -2103 1032 -1991 1038
rect -1925 1072 -1813 1078
rect -1925 1038 -1913 1072
rect -1825 1038 -1813 1072
rect -1925 1032 -1813 1038
rect -1747 1072 -1635 1078
rect -1747 1038 -1735 1072
rect -1647 1038 -1635 1072
rect -1747 1032 -1635 1038
rect -1569 1072 -1457 1078
rect -1569 1038 -1557 1072
rect -1469 1038 -1457 1072
rect -1569 1032 -1457 1038
rect -1391 1072 -1279 1078
rect -1391 1038 -1379 1072
rect -1291 1038 -1279 1072
rect -1391 1032 -1279 1038
rect -1213 1072 -1101 1078
rect -1213 1038 -1201 1072
rect -1113 1038 -1101 1072
rect -1213 1032 -1101 1038
rect -1035 1072 -923 1078
rect -1035 1038 -1023 1072
rect -935 1038 -923 1072
rect -1035 1032 -923 1038
rect -857 1072 -745 1078
rect -857 1038 -845 1072
rect -757 1038 -745 1072
rect -857 1032 -745 1038
rect -679 1072 -567 1078
rect -679 1038 -667 1072
rect -579 1038 -567 1072
rect -679 1032 -567 1038
rect -501 1072 -389 1078
rect -501 1038 -489 1072
rect -401 1038 -389 1072
rect -501 1032 -389 1038
rect -323 1072 -211 1078
rect -323 1038 -311 1072
rect -223 1038 -211 1072
rect -323 1032 -211 1038
rect -145 1072 -33 1078
rect -145 1038 -133 1072
rect -45 1038 -33 1072
rect -145 1032 -33 1038
rect 33 1072 145 1078
rect 33 1038 45 1072
rect 133 1038 145 1072
rect 33 1032 145 1038
rect 211 1072 323 1078
rect 211 1038 223 1072
rect 311 1038 323 1072
rect 211 1032 323 1038
rect 389 1072 501 1078
rect 389 1038 401 1072
rect 489 1038 501 1072
rect 389 1032 501 1038
rect 567 1072 679 1078
rect 567 1038 579 1072
rect 667 1038 679 1072
rect 567 1032 679 1038
rect 745 1072 857 1078
rect 745 1038 757 1072
rect 845 1038 857 1072
rect 745 1032 857 1038
rect 923 1072 1035 1078
rect 923 1038 935 1072
rect 1023 1038 1035 1072
rect 923 1032 1035 1038
rect 1101 1072 1213 1078
rect 1101 1038 1113 1072
rect 1201 1038 1213 1072
rect 1101 1032 1213 1038
rect 1279 1072 1391 1078
rect 1279 1038 1291 1072
rect 1379 1038 1391 1072
rect 1279 1032 1391 1038
rect 1457 1072 1569 1078
rect 1457 1038 1469 1072
rect 1557 1038 1569 1072
rect 1457 1032 1569 1038
rect 1635 1072 1747 1078
rect 1635 1038 1647 1072
rect 1735 1038 1747 1072
rect 1635 1032 1747 1038
rect 1813 1072 1925 1078
rect 1813 1038 1825 1072
rect 1913 1038 1925 1072
rect 1813 1032 1925 1038
rect 1991 1072 2103 1078
rect 1991 1038 2003 1072
rect 2091 1038 2103 1072
rect 1991 1032 2103 1038
rect 2169 1072 2281 1078
rect 2169 1038 2181 1072
rect 2269 1038 2281 1072
rect 2169 1032 2281 1038
rect 2347 1072 2459 1078
rect 2347 1038 2359 1072
rect 2447 1038 2459 1072
rect 2347 1032 2459 1038
rect 2525 1072 2637 1078
rect 2525 1038 2537 1072
rect 2625 1038 2637 1072
rect 2525 1032 2637 1038
rect 2703 1072 2815 1078
rect 2703 1038 2715 1072
rect 2803 1038 2815 1072
rect 2703 1032 2815 1038
rect 2881 1072 2993 1078
rect 2881 1038 2893 1072
rect 2981 1038 2993 1072
rect 2881 1032 2993 1038
rect 3059 1072 3171 1078
rect 3059 1038 3071 1072
rect 3159 1038 3171 1072
rect 3059 1032 3171 1038
rect 3237 1072 3349 1078
rect 3237 1038 3249 1072
rect 3337 1038 3349 1072
rect 3237 1032 3349 1038
rect 3415 1072 3527 1078
rect 3415 1038 3427 1072
rect 3515 1038 3527 1072
rect 3415 1032 3527 1038
rect 3593 1072 3705 1078
rect 3593 1038 3605 1072
rect 3693 1038 3705 1072
rect 3593 1032 3705 1038
rect 3771 1072 3883 1078
rect 3771 1038 3783 1072
rect 3871 1038 3883 1072
rect 3771 1032 3883 1038
rect 3949 1072 4061 1078
rect 3949 1038 3961 1072
rect 4049 1038 4061 1072
rect 3949 1032 4061 1038
rect 4127 1072 4239 1078
rect 4127 1038 4139 1072
rect 4227 1038 4239 1072
rect 4127 1032 4239 1038
rect 4305 1072 4417 1078
rect 4305 1038 4317 1072
rect 4405 1038 4417 1072
rect 4305 1032 4417 1038
rect 4483 1072 4595 1078
rect 4483 1038 4495 1072
rect 4583 1038 4595 1072
rect 4483 1032 4595 1038
rect 4661 1072 4773 1078
rect 4661 1038 4673 1072
rect 4761 1038 4773 1072
rect 4661 1032 4773 1038
rect 4839 1072 4951 1078
rect 4839 1038 4851 1072
rect 4939 1038 4951 1072
rect 4839 1032 4951 1038
rect 5017 1072 5129 1078
rect 5017 1038 5029 1072
rect 5117 1038 5129 1072
rect 5017 1032 5129 1038
rect 5195 1072 5307 1078
rect 5195 1038 5207 1072
rect 5295 1038 5307 1072
rect 5195 1032 5307 1038
rect 5373 1072 5485 1078
rect 5373 1038 5385 1072
rect 5473 1038 5485 1072
rect 5373 1032 5485 1038
rect -5541 988 -5495 1000
rect -5541 -988 -5535 988
rect -5501 -988 -5495 988
rect -5541 -1000 -5495 -988
rect -5363 988 -5317 1000
rect -5363 -988 -5357 988
rect -5323 -988 -5317 988
rect -5363 -1000 -5317 -988
rect -5185 988 -5139 1000
rect -5185 -988 -5179 988
rect -5145 -988 -5139 988
rect -5185 -1000 -5139 -988
rect -5007 988 -4961 1000
rect -5007 -988 -5001 988
rect -4967 -988 -4961 988
rect -5007 -1000 -4961 -988
rect -4829 988 -4783 1000
rect -4829 -988 -4823 988
rect -4789 -988 -4783 988
rect -4829 -1000 -4783 -988
rect -4651 988 -4605 1000
rect -4651 -988 -4645 988
rect -4611 -988 -4605 988
rect -4651 -1000 -4605 -988
rect -4473 988 -4427 1000
rect -4473 -988 -4467 988
rect -4433 -988 -4427 988
rect -4473 -1000 -4427 -988
rect -4295 988 -4249 1000
rect -4295 -988 -4289 988
rect -4255 -988 -4249 988
rect -4295 -1000 -4249 -988
rect -4117 988 -4071 1000
rect -4117 -988 -4111 988
rect -4077 -988 -4071 988
rect -4117 -1000 -4071 -988
rect -3939 988 -3893 1000
rect -3939 -988 -3933 988
rect -3899 -988 -3893 988
rect -3939 -1000 -3893 -988
rect -3761 988 -3715 1000
rect -3761 -988 -3755 988
rect -3721 -988 -3715 988
rect -3761 -1000 -3715 -988
rect -3583 988 -3537 1000
rect -3583 -988 -3577 988
rect -3543 -988 -3537 988
rect -3583 -1000 -3537 -988
rect -3405 988 -3359 1000
rect -3405 -988 -3399 988
rect -3365 -988 -3359 988
rect -3405 -1000 -3359 -988
rect -3227 988 -3181 1000
rect -3227 -988 -3221 988
rect -3187 -988 -3181 988
rect -3227 -1000 -3181 -988
rect -3049 988 -3003 1000
rect -3049 -988 -3043 988
rect -3009 -988 -3003 988
rect -3049 -1000 -3003 -988
rect -2871 988 -2825 1000
rect -2871 -988 -2865 988
rect -2831 -988 -2825 988
rect -2871 -1000 -2825 -988
rect -2693 988 -2647 1000
rect -2693 -988 -2687 988
rect -2653 -988 -2647 988
rect -2693 -1000 -2647 -988
rect -2515 988 -2469 1000
rect -2515 -988 -2509 988
rect -2475 -988 -2469 988
rect -2515 -1000 -2469 -988
rect -2337 988 -2291 1000
rect -2337 -988 -2331 988
rect -2297 -988 -2291 988
rect -2337 -1000 -2291 -988
rect -2159 988 -2113 1000
rect -2159 -988 -2153 988
rect -2119 -988 -2113 988
rect -2159 -1000 -2113 -988
rect -1981 988 -1935 1000
rect -1981 -988 -1975 988
rect -1941 -988 -1935 988
rect -1981 -1000 -1935 -988
rect -1803 988 -1757 1000
rect -1803 -988 -1797 988
rect -1763 -988 -1757 988
rect -1803 -1000 -1757 -988
rect -1625 988 -1579 1000
rect -1625 -988 -1619 988
rect -1585 -988 -1579 988
rect -1625 -1000 -1579 -988
rect -1447 988 -1401 1000
rect -1447 -988 -1441 988
rect -1407 -988 -1401 988
rect -1447 -1000 -1401 -988
rect -1269 988 -1223 1000
rect -1269 -988 -1263 988
rect -1229 -988 -1223 988
rect -1269 -1000 -1223 -988
rect -1091 988 -1045 1000
rect -1091 -988 -1085 988
rect -1051 -988 -1045 988
rect -1091 -1000 -1045 -988
rect -913 988 -867 1000
rect -913 -988 -907 988
rect -873 -988 -867 988
rect -913 -1000 -867 -988
rect -735 988 -689 1000
rect -735 -988 -729 988
rect -695 -988 -689 988
rect -735 -1000 -689 -988
rect -557 988 -511 1000
rect -557 -988 -551 988
rect -517 -988 -511 988
rect -557 -1000 -511 -988
rect -379 988 -333 1000
rect -379 -988 -373 988
rect -339 -988 -333 988
rect -379 -1000 -333 -988
rect -201 988 -155 1000
rect -201 -988 -195 988
rect -161 -988 -155 988
rect -201 -1000 -155 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 155 988 201 1000
rect 155 -988 161 988
rect 195 -988 201 988
rect 155 -1000 201 -988
rect 333 988 379 1000
rect 333 -988 339 988
rect 373 -988 379 988
rect 333 -1000 379 -988
rect 511 988 557 1000
rect 511 -988 517 988
rect 551 -988 557 988
rect 511 -1000 557 -988
rect 689 988 735 1000
rect 689 -988 695 988
rect 729 -988 735 988
rect 689 -1000 735 -988
rect 867 988 913 1000
rect 867 -988 873 988
rect 907 -988 913 988
rect 867 -1000 913 -988
rect 1045 988 1091 1000
rect 1045 -988 1051 988
rect 1085 -988 1091 988
rect 1045 -1000 1091 -988
rect 1223 988 1269 1000
rect 1223 -988 1229 988
rect 1263 -988 1269 988
rect 1223 -1000 1269 -988
rect 1401 988 1447 1000
rect 1401 -988 1407 988
rect 1441 -988 1447 988
rect 1401 -1000 1447 -988
rect 1579 988 1625 1000
rect 1579 -988 1585 988
rect 1619 -988 1625 988
rect 1579 -1000 1625 -988
rect 1757 988 1803 1000
rect 1757 -988 1763 988
rect 1797 -988 1803 988
rect 1757 -1000 1803 -988
rect 1935 988 1981 1000
rect 1935 -988 1941 988
rect 1975 -988 1981 988
rect 1935 -1000 1981 -988
rect 2113 988 2159 1000
rect 2113 -988 2119 988
rect 2153 -988 2159 988
rect 2113 -1000 2159 -988
rect 2291 988 2337 1000
rect 2291 -988 2297 988
rect 2331 -988 2337 988
rect 2291 -1000 2337 -988
rect 2469 988 2515 1000
rect 2469 -988 2475 988
rect 2509 -988 2515 988
rect 2469 -1000 2515 -988
rect 2647 988 2693 1000
rect 2647 -988 2653 988
rect 2687 -988 2693 988
rect 2647 -1000 2693 -988
rect 2825 988 2871 1000
rect 2825 -988 2831 988
rect 2865 -988 2871 988
rect 2825 -1000 2871 -988
rect 3003 988 3049 1000
rect 3003 -988 3009 988
rect 3043 -988 3049 988
rect 3003 -1000 3049 -988
rect 3181 988 3227 1000
rect 3181 -988 3187 988
rect 3221 -988 3227 988
rect 3181 -1000 3227 -988
rect 3359 988 3405 1000
rect 3359 -988 3365 988
rect 3399 -988 3405 988
rect 3359 -1000 3405 -988
rect 3537 988 3583 1000
rect 3537 -988 3543 988
rect 3577 -988 3583 988
rect 3537 -1000 3583 -988
rect 3715 988 3761 1000
rect 3715 -988 3721 988
rect 3755 -988 3761 988
rect 3715 -1000 3761 -988
rect 3893 988 3939 1000
rect 3893 -988 3899 988
rect 3933 -988 3939 988
rect 3893 -1000 3939 -988
rect 4071 988 4117 1000
rect 4071 -988 4077 988
rect 4111 -988 4117 988
rect 4071 -1000 4117 -988
rect 4249 988 4295 1000
rect 4249 -988 4255 988
rect 4289 -988 4295 988
rect 4249 -1000 4295 -988
rect 4427 988 4473 1000
rect 4427 -988 4433 988
rect 4467 -988 4473 988
rect 4427 -1000 4473 -988
rect 4605 988 4651 1000
rect 4605 -988 4611 988
rect 4645 -988 4651 988
rect 4605 -1000 4651 -988
rect 4783 988 4829 1000
rect 4783 -988 4789 988
rect 4823 -988 4829 988
rect 4783 -1000 4829 -988
rect 4961 988 5007 1000
rect 4961 -988 4967 988
rect 5001 -988 5007 988
rect 4961 -1000 5007 -988
rect 5139 988 5185 1000
rect 5139 -988 5145 988
rect 5179 -988 5185 988
rect 5139 -1000 5185 -988
rect 5317 988 5363 1000
rect 5317 -988 5323 988
rect 5357 -988 5363 988
rect 5317 -1000 5363 -988
rect 5495 988 5541 1000
rect 5495 -988 5501 988
rect 5535 -988 5541 988
rect 5495 -1000 5541 -988
rect -5485 -1038 -5373 -1032
rect -5485 -1072 -5473 -1038
rect -5385 -1072 -5373 -1038
rect -5485 -1078 -5373 -1072
rect -5307 -1038 -5195 -1032
rect -5307 -1072 -5295 -1038
rect -5207 -1072 -5195 -1038
rect -5307 -1078 -5195 -1072
rect -5129 -1038 -5017 -1032
rect -5129 -1072 -5117 -1038
rect -5029 -1072 -5017 -1038
rect -5129 -1078 -5017 -1072
rect -4951 -1038 -4839 -1032
rect -4951 -1072 -4939 -1038
rect -4851 -1072 -4839 -1038
rect -4951 -1078 -4839 -1072
rect -4773 -1038 -4661 -1032
rect -4773 -1072 -4761 -1038
rect -4673 -1072 -4661 -1038
rect -4773 -1078 -4661 -1072
rect -4595 -1038 -4483 -1032
rect -4595 -1072 -4583 -1038
rect -4495 -1072 -4483 -1038
rect -4595 -1078 -4483 -1072
rect -4417 -1038 -4305 -1032
rect -4417 -1072 -4405 -1038
rect -4317 -1072 -4305 -1038
rect -4417 -1078 -4305 -1072
rect -4239 -1038 -4127 -1032
rect -4239 -1072 -4227 -1038
rect -4139 -1072 -4127 -1038
rect -4239 -1078 -4127 -1072
rect -4061 -1038 -3949 -1032
rect -4061 -1072 -4049 -1038
rect -3961 -1072 -3949 -1038
rect -4061 -1078 -3949 -1072
rect -3883 -1038 -3771 -1032
rect -3883 -1072 -3871 -1038
rect -3783 -1072 -3771 -1038
rect -3883 -1078 -3771 -1072
rect -3705 -1038 -3593 -1032
rect -3705 -1072 -3693 -1038
rect -3605 -1072 -3593 -1038
rect -3705 -1078 -3593 -1072
rect -3527 -1038 -3415 -1032
rect -3527 -1072 -3515 -1038
rect -3427 -1072 -3415 -1038
rect -3527 -1078 -3415 -1072
rect -3349 -1038 -3237 -1032
rect -3349 -1072 -3337 -1038
rect -3249 -1072 -3237 -1038
rect -3349 -1078 -3237 -1072
rect -3171 -1038 -3059 -1032
rect -3171 -1072 -3159 -1038
rect -3071 -1072 -3059 -1038
rect -3171 -1078 -3059 -1072
rect -2993 -1038 -2881 -1032
rect -2993 -1072 -2981 -1038
rect -2893 -1072 -2881 -1038
rect -2993 -1078 -2881 -1072
rect -2815 -1038 -2703 -1032
rect -2815 -1072 -2803 -1038
rect -2715 -1072 -2703 -1038
rect -2815 -1078 -2703 -1072
rect -2637 -1038 -2525 -1032
rect -2637 -1072 -2625 -1038
rect -2537 -1072 -2525 -1038
rect -2637 -1078 -2525 -1072
rect -2459 -1038 -2347 -1032
rect -2459 -1072 -2447 -1038
rect -2359 -1072 -2347 -1038
rect -2459 -1078 -2347 -1072
rect -2281 -1038 -2169 -1032
rect -2281 -1072 -2269 -1038
rect -2181 -1072 -2169 -1038
rect -2281 -1078 -2169 -1072
rect -2103 -1038 -1991 -1032
rect -2103 -1072 -2091 -1038
rect -2003 -1072 -1991 -1038
rect -2103 -1078 -1991 -1072
rect -1925 -1038 -1813 -1032
rect -1925 -1072 -1913 -1038
rect -1825 -1072 -1813 -1038
rect -1925 -1078 -1813 -1072
rect -1747 -1038 -1635 -1032
rect -1747 -1072 -1735 -1038
rect -1647 -1072 -1635 -1038
rect -1747 -1078 -1635 -1072
rect -1569 -1038 -1457 -1032
rect -1569 -1072 -1557 -1038
rect -1469 -1072 -1457 -1038
rect -1569 -1078 -1457 -1072
rect -1391 -1038 -1279 -1032
rect -1391 -1072 -1379 -1038
rect -1291 -1072 -1279 -1038
rect -1391 -1078 -1279 -1072
rect -1213 -1038 -1101 -1032
rect -1213 -1072 -1201 -1038
rect -1113 -1072 -1101 -1038
rect -1213 -1078 -1101 -1072
rect -1035 -1038 -923 -1032
rect -1035 -1072 -1023 -1038
rect -935 -1072 -923 -1038
rect -1035 -1078 -923 -1072
rect -857 -1038 -745 -1032
rect -857 -1072 -845 -1038
rect -757 -1072 -745 -1038
rect -857 -1078 -745 -1072
rect -679 -1038 -567 -1032
rect -679 -1072 -667 -1038
rect -579 -1072 -567 -1038
rect -679 -1078 -567 -1072
rect -501 -1038 -389 -1032
rect -501 -1072 -489 -1038
rect -401 -1072 -389 -1038
rect -501 -1078 -389 -1072
rect -323 -1038 -211 -1032
rect -323 -1072 -311 -1038
rect -223 -1072 -211 -1038
rect -323 -1078 -211 -1072
rect -145 -1038 -33 -1032
rect -145 -1072 -133 -1038
rect -45 -1072 -33 -1038
rect -145 -1078 -33 -1072
rect 33 -1038 145 -1032
rect 33 -1072 45 -1038
rect 133 -1072 145 -1038
rect 33 -1078 145 -1072
rect 211 -1038 323 -1032
rect 211 -1072 223 -1038
rect 311 -1072 323 -1038
rect 211 -1078 323 -1072
rect 389 -1038 501 -1032
rect 389 -1072 401 -1038
rect 489 -1072 501 -1038
rect 389 -1078 501 -1072
rect 567 -1038 679 -1032
rect 567 -1072 579 -1038
rect 667 -1072 679 -1038
rect 567 -1078 679 -1072
rect 745 -1038 857 -1032
rect 745 -1072 757 -1038
rect 845 -1072 857 -1038
rect 745 -1078 857 -1072
rect 923 -1038 1035 -1032
rect 923 -1072 935 -1038
rect 1023 -1072 1035 -1038
rect 923 -1078 1035 -1072
rect 1101 -1038 1213 -1032
rect 1101 -1072 1113 -1038
rect 1201 -1072 1213 -1038
rect 1101 -1078 1213 -1072
rect 1279 -1038 1391 -1032
rect 1279 -1072 1291 -1038
rect 1379 -1072 1391 -1038
rect 1279 -1078 1391 -1072
rect 1457 -1038 1569 -1032
rect 1457 -1072 1469 -1038
rect 1557 -1072 1569 -1038
rect 1457 -1078 1569 -1072
rect 1635 -1038 1747 -1032
rect 1635 -1072 1647 -1038
rect 1735 -1072 1747 -1038
rect 1635 -1078 1747 -1072
rect 1813 -1038 1925 -1032
rect 1813 -1072 1825 -1038
rect 1913 -1072 1925 -1038
rect 1813 -1078 1925 -1072
rect 1991 -1038 2103 -1032
rect 1991 -1072 2003 -1038
rect 2091 -1072 2103 -1038
rect 1991 -1078 2103 -1072
rect 2169 -1038 2281 -1032
rect 2169 -1072 2181 -1038
rect 2269 -1072 2281 -1038
rect 2169 -1078 2281 -1072
rect 2347 -1038 2459 -1032
rect 2347 -1072 2359 -1038
rect 2447 -1072 2459 -1038
rect 2347 -1078 2459 -1072
rect 2525 -1038 2637 -1032
rect 2525 -1072 2537 -1038
rect 2625 -1072 2637 -1038
rect 2525 -1078 2637 -1072
rect 2703 -1038 2815 -1032
rect 2703 -1072 2715 -1038
rect 2803 -1072 2815 -1038
rect 2703 -1078 2815 -1072
rect 2881 -1038 2993 -1032
rect 2881 -1072 2893 -1038
rect 2981 -1072 2993 -1038
rect 2881 -1078 2993 -1072
rect 3059 -1038 3171 -1032
rect 3059 -1072 3071 -1038
rect 3159 -1072 3171 -1038
rect 3059 -1078 3171 -1072
rect 3237 -1038 3349 -1032
rect 3237 -1072 3249 -1038
rect 3337 -1072 3349 -1038
rect 3237 -1078 3349 -1072
rect 3415 -1038 3527 -1032
rect 3415 -1072 3427 -1038
rect 3515 -1072 3527 -1038
rect 3415 -1078 3527 -1072
rect 3593 -1038 3705 -1032
rect 3593 -1072 3605 -1038
rect 3693 -1072 3705 -1038
rect 3593 -1078 3705 -1072
rect 3771 -1038 3883 -1032
rect 3771 -1072 3783 -1038
rect 3871 -1072 3883 -1038
rect 3771 -1078 3883 -1072
rect 3949 -1038 4061 -1032
rect 3949 -1072 3961 -1038
rect 4049 -1072 4061 -1038
rect 3949 -1078 4061 -1072
rect 4127 -1038 4239 -1032
rect 4127 -1072 4139 -1038
rect 4227 -1072 4239 -1038
rect 4127 -1078 4239 -1072
rect 4305 -1038 4417 -1032
rect 4305 -1072 4317 -1038
rect 4405 -1072 4417 -1038
rect 4305 -1078 4417 -1072
rect 4483 -1038 4595 -1032
rect 4483 -1072 4495 -1038
rect 4583 -1072 4595 -1038
rect 4483 -1078 4595 -1072
rect 4661 -1038 4773 -1032
rect 4661 -1072 4673 -1038
rect 4761 -1072 4773 -1038
rect 4661 -1078 4773 -1072
rect 4839 -1038 4951 -1032
rect 4839 -1072 4851 -1038
rect 4939 -1072 4951 -1038
rect 4839 -1078 4951 -1072
rect 5017 -1038 5129 -1032
rect 5017 -1072 5029 -1038
rect 5117 -1072 5129 -1038
rect 5017 -1078 5129 -1072
rect 5195 -1038 5307 -1032
rect 5195 -1072 5207 -1038
rect 5295 -1072 5307 -1038
rect 5195 -1078 5307 -1072
rect 5373 -1038 5485 -1032
rect 5373 -1072 5385 -1038
rect 5473 -1072 5485 -1038
rect 5373 -1078 5485 -1072
<< properties >>
string FIXED_BBOX -5632 -1157 5632 1157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 0.6 m 1 nf 62 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
