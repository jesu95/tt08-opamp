magic
tech sky130A
magscale 1 2
timestamp 1723396918
<< nwell >>
rect 2786 30924 5024 38338
rect 4556 8432 6794 15740
<< pwell >>
rect 20894 40044 23264 40102
rect 20898 39806 23268 39864
rect 20892 37686 23262 37744
rect 20910 37448 23280 37506
rect 20906 37214 23276 37272
rect 20932 36978 23302 37036
rect 20920 36740 23290 36798
rect 20892 36502 23262 36560
rect 20884 36270 23254 36328
rect 20920 36034 23290 36092
rect 20912 35796 23282 35854
rect 20900 35562 23270 35620
rect 20952 35326 23322 35384
rect 20934 35090 23304 35148
rect 21004 34618 23374 34676
rect 20942 34382 23312 34440
rect 20880 34144 23250 34202
rect 20900 33908 23270 33966
rect 20938 33674 23308 33732
rect 20940 33436 23310 33494
rect 20900 33200 23270 33258
rect 20894 32966 23264 33024
rect 20950 32730 23320 32788
rect 20936 32492 23306 32550
rect 20974 32256 23344 32314
rect 20948 32020 23318 32078
rect 20928 31782 23298 31840
rect 20900 31548 23270 31606
rect 20908 31314 23278 31372
rect 20900 31078 23270 31136
rect 20884 30840 23254 30898
rect 20960 30604 23330 30662
rect 21112 30368 23482 30426
rect 21062 30132 23432 30190
rect 23068 2840 23170 25042
<< pdiff >>
rect 4782 15298 6570 15352
rect 4782 14354 6570 14408
rect 4782 11286 6570 11340
<< locali >>
rect 23260 44452 27492 44454
rect 1996 38266 4954 44450
rect 20460 43860 27492 44452
rect 20460 43240 23738 43860
rect 27086 43240 27492 43860
rect 20460 40588 27492 43240
rect 20460 40520 25116 40588
rect 1996 30994 2860 38266
rect 1996 30458 4968 30994
rect 1996 29890 4966 30458
rect 1996 3110 2784 29890
rect 3772 22968 4966 29890
rect 23180 29710 25116 40520
rect 20460 25840 25116 29710
rect 20460 25440 20524 25840
rect 20670 25440 25116 25840
rect 20460 25280 25116 25440
rect 3772 21812 6198 22968
rect 3772 21412 5598 21812
rect 5998 21412 6198 21812
rect 3772 15776 6198 21412
rect 3772 7568 4628 15776
rect 3772 3110 6194 7568
rect 1996 2802 6194 3110
rect 23180 2804 25116 25280
rect 1996 1000 19742 2802
rect 20864 2770 23210 2804
rect 23212 2770 25116 2804
rect 20864 2734 25116 2770
rect 25640 2734 27492 40588
rect 20864 1000 27492 2734
<< viali >>
rect 23738 43240 27086 43860
rect 2784 3110 3772 29890
rect 20524 25440 20670 25840
rect 5598 21412 5998 21812
rect 19722 21594 19760 21684
rect 25116 2734 25640 40588
<< metal1 >>
rect 23726 43860 27098 43866
rect 23726 43240 23738 43860
rect 27086 43240 27098 43860
rect 23726 43234 27098 43240
rect 25110 40588 25646 40600
rect 4838 38302 5194 38304
rect 3018 38204 4792 38214
rect 2874 30924 2972 38182
rect 3018 38128 4792 38138
rect 3012 38080 4800 38090
rect 3012 38016 4800 38026
rect 3018 37968 4792 37978
rect 3018 37892 4792 37902
rect 3012 37844 4800 37854
rect 3012 37780 4800 37790
rect 3018 37732 4792 37742
rect 3018 37656 4792 37666
rect 3012 37608 4800 37618
rect 3012 37544 4800 37554
rect 3018 37496 4792 37506
rect 3018 37420 4792 37430
rect 3012 37372 4800 37382
rect 3012 37308 4800 37318
rect 3018 37260 4792 37270
rect 3018 37184 4792 37194
rect 3012 37136 4800 37146
rect 3012 37072 4800 37082
rect 3018 37024 4792 37034
rect 3018 36948 4792 36958
rect 3012 36900 4800 36910
rect 3012 36836 4800 36846
rect 3018 36788 4792 36798
rect 3018 36712 4792 36722
rect 3012 36664 4800 36674
rect 3012 36600 4800 36610
rect 3018 36552 4792 36562
rect 3018 36476 4792 36486
rect 3012 36428 4800 36438
rect 3012 36364 4800 36374
rect 3018 36316 4792 36326
rect 3018 36240 4792 36250
rect 3012 36192 4800 36202
rect 3012 36128 4800 36138
rect 3018 36080 4792 36090
rect 3018 36004 4792 36014
rect 3012 35956 4800 35966
rect 3012 35892 4800 35902
rect 3018 35844 4792 35854
rect 3018 35768 4792 35778
rect 3012 35720 4800 35730
rect 3012 35656 4800 35666
rect 3018 35608 4792 35618
rect 3018 35532 4792 35542
rect 3012 35484 4800 35494
rect 3012 35420 4800 35430
rect 3018 35372 4792 35382
rect 3018 35296 4792 35306
rect 3012 35248 4800 35258
rect 3012 35184 4800 35194
rect 3018 35136 4792 35146
rect 3018 35060 4792 35070
rect 3012 35012 4800 35022
rect 3012 34948 4800 34958
rect 3018 34900 4792 34910
rect 3018 34824 4792 34834
rect 3012 34776 4800 34786
rect 3012 34712 4800 34722
rect 3018 34664 4792 34674
rect 3018 34588 4792 34598
rect 3012 34540 4800 34550
rect 3012 34476 4800 34486
rect 3018 34428 4792 34438
rect 3018 34352 4792 34362
rect 3012 34304 4800 34314
rect 3012 34240 4800 34250
rect 3018 34192 4792 34202
rect 3018 34116 4792 34126
rect 3012 34068 4800 34078
rect 3012 34004 4800 34014
rect 3018 33956 4792 33966
rect 3018 33880 4792 33890
rect 3012 33832 4800 33842
rect 3012 33768 4800 33778
rect 3018 33720 4792 33730
rect 3018 33644 4792 33654
rect 3012 33596 4800 33606
rect 3012 33532 4800 33542
rect 3018 33484 4792 33494
rect 3018 33408 4792 33418
rect 3012 33360 4800 33370
rect 3012 33296 4800 33306
rect 3018 33248 4792 33258
rect 3018 33172 4792 33182
rect 3012 33124 4800 33134
rect 3012 33060 4800 33070
rect 3018 33012 4792 33022
rect 3018 32936 4792 32946
rect 3012 32888 4800 32898
rect 3012 32824 4800 32834
rect 3018 32776 4792 32786
rect 3018 32700 4792 32710
rect 3012 32652 4800 32662
rect 3012 32588 4800 32598
rect 3018 32540 4792 32550
rect 3018 32464 4792 32474
rect 3012 32416 4800 32426
rect 3012 32352 4800 32362
rect 3018 32304 4792 32314
rect 3018 32228 4792 32238
rect 3012 32180 4800 32190
rect 3012 32116 4800 32126
rect 3018 32068 4792 32078
rect 3018 31992 4792 32002
rect 3012 31944 4800 31954
rect 3012 31880 4800 31890
rect 3016 31832 4790 31842
rect 3016 31756 4790 31766
rect 3012 31708 4800 31718
rect 3012 31644 4800 31654
rect 3018 31596 4792 31606
rect 3018 31520 4792 31530
rect 3012 31472 4800 31482
rect 3012 31408 4800 31418
rect 3018 31360 4792 31370
rect 3018 31284 4792 31294
rect 3012 31236 4800 31246
rect 3012 31172 4800 31182
rect 3018 31120 4792 31130
rect 3018 31050 4792 31060
rect 2778 29890 3778 29902
rect 2774 3110 2784 29890
rect 3772 3110 3782 29890
rect 4836 20606 5194 38302
rect 20520 29640 20612 40470
rect 20656 40460 23026 40470
rect 20656 40386 23026 40396
rect 20658 40338 23028 40348
rect 20658 40270 23028 40280
rect 20656 40224 23026 40234
rect 20656 40150 23026 40160
rect 20656 40104 23026 40114
rect 20656 40036 23026 40046
rect 20654 39988 23024 39998
rect 20654 39914 23024 39924
rect 20658 39864 23028 39874
rect 20658 39796 23028 39806
rect 20654 39752 23024 39762
rect 20654 39678 23024 39688
rect 20656 39632 23026 39642
rect 20656 39564 23026 39574
rect 20656 39516 23026 39526
rect 20656 39442 23026 39452
rect 20656 39394 23026 39404
rect 20656 39326 23026 39336
rect 20654 39278 23024 39288
rect 20654 39204 23024 39214
rect 20656 39160 23026 39170
rect 20656 39092 23026 39102
rect 20656 39042 23026 39052
rect 20656 38968 23026 38978
rect 20656 38924 23026 38934
rect 20656 38856 23026 38866
rect 20654 38810 23024 38820
rect 20654 38736 23024 38746
rect 20658 38686 23028 38696
rect 20658 38618 23028 38628
rect 20656 38570 23026 38580
rect 20656 38496 23026 38506
rect 20656 38450 23026 38460
rect 20656 38382 23026 38392
rect 20654 38334 23024 38344
rect 20654 38260 23024 38270
rect 20656 38214 23026 38224
rect 20656 38146 23026 38156
rect 20654 38098 23024 38108
rect 20654 38024 23024 38034
rect 20656 37978 23026 37988
rect 20656 37910 23026 37920
rect 20656 37862 23026 37872
rect 20656 37788 23026 37798
rect 20658 37744 23028 37754
rect 20658 37676 23028 37686
rect 20656 37626 23026 37636
rect 20656 37552 23026 37562
rect 20656 37506 23026 37516
rect 20656 37438 23026 37448
rect 20656 37390 23026 37400
rect 20656 37316 23026 37326
rect 20658 37268 23028 37278
rect 20658 37200 23028 37210
rect 20654 37156 23024 37166
rect 20654 37082 23024 37092
rect 20658 37034 23028 37044
rect 20658 36966 23028 36976
rect 20658 36920 23028 36930
rect 20658 36846 23028 36856
rect 20658 36798 23028 36808
rect 20658 36730 23028 36740
rect 20656 36682 23026 36692
rect 20656 36608 23026 36618
rect 20656 36562 23026 36572
rect 20656 36494 23026 36504
rect 20658 36446 23028 36456
rect 20658 36372 23028 36382
rect 20658 36326 23028 36336
rect 20658 36258 23028 36268
rect 20658 36210 23028 36220
rect 20658 36136 23028 36146
rect 20656 36090 23026 36100
rect 20656 36022 23026 36032
rect 20658 35976 23028 35986
rect 20658 35902 23028 35912
rect 20656 35856 23026 35866
rect 20656 35788 23026 35798
rect 20654 35738 23024 35748
rect 20654 35664 23024 35674
rect 20658 35620 23028 35630
rect 20658 35552 23028 35562
rect 20654 35500 23024 35510
rect 20654 35426 23024 35436
rect 20656 35384 23026 35394
rect 20656 35316 23026 35326
rect 20656 35266 23026 35276
rect 20656 35192 23026 35202
rect 20656 35148 23026 35158
rect 20656 35080 23026 35090
rect 20656 35030 23026 35040
rect 20656 34956 23026 34966
rect 20656 34910 23026 34920
rect 20656 34842 23026 34852
rect 20658 34794 23028 34804
rect 20658 34720 23028 34730
rect 20658 34674 23028 34684
rect 20658 34606 23028 34616
rect 20654 34560 23024 34570
rect 20654 34486 23024 34496
rect 20660 34438 23030 34448
rect 20660 34370 23030 34380
rect 20654 34322 23024 34332
rect 20654 34248 23024 34258
rect 20658 34202 23028 34212
rect 20658 34134 23028 34144
rect 20656 34088 23026 34098
rect 20656 34014 23026 34024
rect 20656 33964 23026 33974
rect 20656 33896 23026 33906
rect 20656 33850 23026 33860
rect 20656 33776 23026 33786
rect 20656 33732 23026 33742
rect 20656 33664 23026 33674
rect 20656 33614 23026 33624
rect 20656 33540 23026 33550
rect 20656 33494 23026 33504
rect 20656 33426 23026 33436
rect 20656 33380 23026 33390
rect 20656 33306 23026 33316
rect 20658 33260 23028 33270
rect 20658 33192 23028 33202
rect 20656 33144 23026 33154
rect 20656 33070 23026 33080
rect 20658 33022 23028 33032
rect 20658 32954 23028 32964
rect 20656 32906 23026 32916
rect 20656 32832 23026 32842
rect 20656 32788 23026 32798
rect 20656 32720 23026 32730
rect 20658 32672 23028 32682
rect 20658 32598 23028 32608
rect 20656 32552 23026 32562
rect 20656 32484 23026 32494
rect 20658 32438 23028 32448
rect 20658 32364 23028 32374
rect 20656 32314 23026 32324
rect 20656 32246 23026 32256
rect 20656 32198 23026 32208
rect 20656 32124 23026 32134
rect 20656 32078 23026 32088
rect 20656 32010 23026 32020
rect 20656 31964 23026 31974
rect 20656 31890 23026 31900
rect 20658 31840 23028 31850
rect 20658 31772 23028 31782
rect 20656 31726 23026 31736
rect 20656 31652 23026 31662
rect 20658 31606 23028 31616
rect 20658 31538 23028 31548
rect 20656 31492 23026 31502
rect 20656 31418 23026 31428
rect 20658 31372 23028 31382
rect 20658 31304 23028 31314
rect 20656 31256 23026 31266
rect 20656 31182 23026 31192
rect 20656 31134 23026 31144
rect 20656 31066 23026 31076
rect 20654 31020 23024 31030
rect 20654 30946 23024 30956
rect 20656 30900 23026 30910
rect 20656 30832 23026 30842
rect 20656 30782 23026 30792
rect 20656 30708 23026 30718
rect 20656 30662 23026 30672
rect 20656 30594 23026 30604
rect 20656 30546 23026 30556
rect 20656 30472 23026 30482
rect 20656 30426 23026 30436
rect 20656 30358 23026 30368
rect 20656 30312 23026 30322
rect 20656 30238 23026 30248
rect 20658 30188 23028 30198
rect 20658 30120 23028 30130
rect 20656 30074 23026 30084
rect 20656 30000 23026 30010
rect 20658 29954 23028 29964
rect 20658 29886 23028 29896
rect 20658 29840 23028 29850
rect 20658 29766 23028 29776
rect 23070 29738 23172 40494
rect 20476 27440 20676 29640
rect 19788 27244 20676 27440
rect 19788 22772 19996 27244
rect 18468 22294 18478 22684
rect 18982 22648 18992 22684
rect 19788 22660 19814 22772
rect 19974 22660 19996 22772
rect 19788 22648 19996 22660
rect 20492 25840 20702 26040
rect 20492 25440 20524 25840
rect 20670 25440 20702 25840
rect 18982 22294 18992 22330
rect 5544 21812 17754 21930
rect 5544 21412 5598 21812
rect 5998 21412 17754 21812
rect 18522 21688 18922 22294
rect 20492 21818 20702 25440
rect 19722 21696 20702 21818
rect 19716 21684 20702 21696
rect 5544 21340 17754 21412
rect 18522 21154 18924 21596
rect 19716 21594 19722 21684
rect 19760 21594 20702 21684
rect 19716 21582 20702 21594
rect 19722 21534 20702 21582
rect 20904 25168 21006 25240
rect 21052 25226 23024 25236
rect 19722 21466 20700 21534
rect 19738 21464 19774 21466
rect 18522 21144 19994 21154
rect 18522 21030 19810 21144
rect 19970 21030 19994 21144
rect 18522 21020 19994 21030
rect 9172 20730 11542 20740
rect 9172 20656 11542 20666
rect 4836 20112 6996 20606
rect 9174 20556 11542 20566
rect 9172 20486 9174 20556
rect 9174 20476 11542 20486
rect 9172 20374 11542 20384
rect 9172 20300 11542 20310
rect 9172 20200 11540 20210
rect 9172 20120 11540 20130
rect 4838 20110 5194 20112
rect 6500 16040 6994 20112
rect 9172 20018 11542 20028
rect 9172 19944 11542 19954
rect 9172 19844 11540 19854
rect 9172 19764 11540 19774
rect 9172 19662 11542 19672
rect 9172 19588 11542 19598
rect 9172 19490 11540 19500
rect 9172 19410 11540 19420
rect 9172 19308 11542 19318
rect 9172 19234 11542 19244
rect 9172 19132 11540 19142
rect 9172 19052 11540 19062
rect 9172 18950 11542 18960
rect 9172 18876 11542 18886
rect 9172 18776 11540 18786
rect 9172 18696 11540 18706
rect 9172 18594 11542 18604
rect 9172 18520 11542 18530
rect 9172 18420 11540 18430
rect 9172 18340 11540 18350
rect 9172 18238 11542 18248
rect 9172 18164 11542 18174
rect 9172 18064 11540 18074
rect 9172 17984 11540 17994
rect 9172 17882 11542 17892
rect 9172 17808 11542 17818
rect 9172 17708 11540 17718
rect 9172 17628 11540 17638
rect 9172 17528 11542 17538
rect 9172 17454 11542 17464
rect 9172 17350 11540 17360
rect 9172 17270 11540 17280
rect 9172 17172 11542 17182
rect 9172 17098 11542 17108
rect 9172 16996 11540 17006
rect 9172 16916 11540 16926
rect 9172 16816 11542 16826
rect 9172 16742 11542 16752
rect 9172 16640 11540 16650
rect 9172 16560 11540 16570
rect 9172 16462 11542 16472
rect 9172 16388 11542 16398
rect 9172 16286 11540 16296
rect 9172 16206 11540 16216
rect 9172 16102 11542 16112
rect 6610 15740 6876 16040
rect 9172 16028 11542 16038
rect 9172 15928 11540 15938
rect 9172 15848 11540 15858
rect 4644 7632 4742 15740
rect 4780 15710 6568 15720
rect 4780 15638 6568 15648
rect 4782 15588 6570 15598
rect 4782 15524 6570 15534
rect 4780 15474 6568 15484
rect 4780 15402 6568 15412
rect 4782 15352 6570 15362
rect 4782 15288 6570 15298
rect 4780 15238 6568 15248
rect 4780 15166 6568 15176
rect 4782 15116 6570 15126
rect 4782 15052 6570 15062
rect 4780 15002 6568 15012
rect 4780 14930 6568 14940
rect 4782 14880 6570 14890
rect 4782 14816 6570 14826
rect 4780 14766 6568 14776
rect 4780 14694 6568 14704
rect 4782 14644 6570 14654
rect 4782 14580 6570 14590
rect 4780 14530 6568 14540
rect 4780 14458 6568 14468
rect 4782 14408 6570 14418
rect 4782 14344 6570 14354
rect 4780 14294 6568 14304
rect 4780 14222 6568 14232
rect 4780 14172 6568 14182
rect 4780 14108 6568 14118
rect 4778 14058 6566 14068
rect 6566 13996 6568 14058
rect 4778 13986 6566 13996
rect 4780 13936 6568 13946
rect 4780 13872 6568 13882
rect 4780 13822 6568 13832
rect 4780 13750 6568 13760
rect 4782 13700 6570 13710
rect 4782 13636 6570 13646
rect 4780 13586 6568 13596
rect 4780 13514 6568 13524
rect 4782 13464 6570 13474
rect 4782 13400 6570 13410
rect 4780 13350 6568 13360
rect 4780 13278 6568 13288
rect 4782 13228 6570 13238
rect 4782 13164 6570 13174
rect 4780 13114 6568 13124
rect 4780 13042 6568 13052
rect 4782 12992 6570 13002
rect 4782 12928 6570 12938
rect 4780 12878 6568 12888
rect 4780 12806 6568 12816
rect 4782 12756 6570 12766
rect 4782 12692 6570 12702
rect 4778 12642 6566 12652
rect 6566 12580 6568 12642
rect 4778 12570 6566 12580
rect 4782 12520 6570 12530
rect 4782 12456 6570 12466
rect 4780 12406 6568 12416
rect 4780 12334 6568 12344
rect 4782 12284 6570 12294
rect 4782 12220 6570 12230
rect 4780 12170 6568 12180
rect 4780 12098 6568 12108
rect 4782 12048 6570 12058
rect 4782 11984 6570 11994
rect 4780 11934 6568 11944
rect 4780 11862 6568 11872
rect 4782 11812 6570 11822
rect 4782 11748 6570 11758
rect 4778 11698 6566 11708
rect 6566 11636 6568 11698
rect 4778 11626 6566 11636
rect 4782 11576 6570 11586
rect 4782 11512 6570 11522
rect 4778 11462 6566 11472
rect 6566 11400 6568 11462
rect 4778 11390 6566 11400
rect 4782 11340 6570 11350
rect 4782 11276 6570 11286
rect 4780 11226 6568 11236
rect 4780 11154 6568 11164
rect 4782 11104 6570 11114
rect 4782 11040 6570 11050
rect 4780 10990 6568 11000
rect 4780 10918 6568 10928
rect 4782 10868 6570 10878
rect 4782 10804 6570 10814
rect 4780 10754 6568 10764
rect 4780 10682 6568 10692
rect 4782 10632 6570 10642
rect 4782 10568 6570 10578
rect 4780 10518 6568 10528
rect 4780 10446 6568 10456
rect 4782 10396 6570 10406
rect 4782 10332 6570 10342
rect 4778 10282 6566 10292
rect 6566 10220 6568 10282
rect 4778 10210 6566 10220
rect 4782 10160 6570 10170
rect 4782 10096 6570 10106
rect 4778 10046 6566 10056
rect 6566 9984 6568 10046
rect 4778 9974 6566 9984
rect 4782 9924 6570 9934
rect 4782 9860 6570 9870
rect 4780 9810 6568 9820
rect 4780 9738 6568 9748
rect 4782 9688 6570 9698
rect 4782 9624 6570 9634
rect 4778 9574 6566 9584
rect 6566 9512 6568 9574
rect 4778 9502 6566 9512
rect 4782 9452 6570 9462
rect 4780 9398 4782 9452
rect 4782 9388 6570 9398
rect 4780 9338 6568 9348
rect 4780 9266 6568 9276
rect 4780 9216 6568 9226
rect 4780 9152 6568 9162
rect 4778 9102 6566 9110
rect 4778 9100 6568 9102
rect 6566 9038 6568 9100
rect 4778 9028 6566 9038
rect 4780 8980 6568 8990
rect 4780 8916 6568 8926
rect 4778 8868 6566 8876
rect 4778 8866 6568 8868
rect 6566 8804 6568 8866
rect 4778 8794 6566 8804
rect 4780 8744 6568 8754
rect 4780 8680 6568 8690
rect 4780 8630 6568 8640
rect 4780 8558 6568 8568
rect 6608 8398 6876 15740
rect 9172 15746 11542 15756
rect 9172 15672 11542 15682
rect 9172 15572 11540 15582
rect 9172 15492 11540 15502
rect 9172 15392 11542 15402
rect 9172 15318 11542 15328
rect 9172 15216 11540 15226
rect 9172 15136 11540 15146
rect 9172 15034 11542 15044
rect 9172 14960 11542 14970
rect 9172 14860 11540 14870
rect 9172 14780 11540 14790
rect 9172 14680 11542 14690
rect 9172 14606 11542 14616
rect 9172 14504 11540 14514
rect 9172 14424 11540 14434
rect 9172 14322 11542 14332
rect 9172 14248 11542 14258
rect 9172 14148 11540 14158
rect 9172 14068 11540 14078
rect 9172 13968 11542 13978
rect 9172 13894 11542 13904
rect 9172 13792 11540 13802
rect 9172 13712 11540 13722
rect 9172 13614 11542 13624
rect 9172 13540 11542 13550
rect 9172 13436 11540 13446
rect 9172 13356 11540 13366
rect 9172 13256 11542 13266
rect 9172 13182 11542 13192
rect 9172 13080 11540 13090
rect 9172 13000 11540 13010
rect 9172 12898 11542 12908
rect 9172 12824 11542 12834
rect 9172 12724 11540 12734
rect 9172 12644 11540 12654
rect 9172 12544 11542 12554
rect 9172 12470 11542 12480
rect 9172 12368 11540 12378
rect 9172 12288 11540 12298
rect 9172 12186 11542 12196
rect 9172 12112 11542 12122
rect 9172 12012 11540 12022
rect 9172 11932 11540 11942
rect 9172 11830 11542 11840
rect 9172 11756 11542 11766
rect 9170 11656 11538 11666
rect 9170 11576 11538 11586
rect 9172 11476 11542 11486
rect 9172 11402 11542 11412
rect 9170 11300 11538 11310
rect 9170 11220 11538 11230
rect 9172 11120 11542 11130
rect 9172 11046 11542 11056
rect 9170 10944 11538 10954
rect 9170 10864 11538 10874
rect 9172 10764 11542 10774
rect 9172 10690 11542 10700
rect 9170 10588 11538 10598
rect 9170 10508 11538 10518
rect 9170 10408 11540 10418
rect 9170 10334 11540 10344
rect 9170 10230 11538 10240
rect 9170 10150 11538 10160
rect 9172 10052 11542 10062
rect 9172 9978 11542 9988
rect 9170 9876 11538 9886
rect 9170 9796 11538 9806
rect 9172 9696 11542 9706
rect 9172 9622 11542 9632
rect 9172 9520 11540 9530
rect 9172 9440 11540 9450
rect 9172 9342 11542 9352
rect 9172 9268 11542 9278
rect 9172 9164 11540 9174
rect 9172 9084 11540 9094
rect 9172 8982 11542 8992
rect 9172 8908 11542 8918
rect 9172 8806 11540 8816
rect 9172 8726 11540 8736
rect 9172 8626 11542 8636
rect 9172 8552 11542 8562
rect 4810 8342 6876 8398
rect 9172 8452 11540 8462
rect 9172 8372 11540 8382
rect 4788 8282 6568 8292
rect 4788 8214 6568 8224
rect 6608 8164 6876 8342
rect 9172 8272 11542 8282
rect 9172 8198 11542 8208
rect 4798 8108 6876 8164
rect 4788 8046 6568 8056
rect 4788 7978 6568 7988
rect 6608 7926 6876 8108
rect 9172 8096 11540 8106
rect 9172 8016 11540 8026
rect 4800 7870 6876 7926
rect 4788 7810 6568 7820
rect 4788 7742 6568 7752
rect 6608 7692 6876 7870
rect 9172 7916 11542 7926
rect 9172 7842 11542 7852
rect 4782 7688 6876 7692
rect 4778 7636 6876 7688
rect 9172 7740 11540 7750
rect 9172 7660 11540 7670
rect 4778 7634 6566 7636
rect 6608 6802 6876 7636
rect 9172 7560 11542 7570
rect 9172 7486 11542 7496
rect 9172 7384 11540 7394
rect 9172 7304 11540 7314
rect 9172 7204 11542 7214
rect 9172 7130 11542 7140
rect 9172 7028 11540 7038
rect 9172 6948 11540 6958
rect 9172 6848 11542 6858
rect 2778 3098 3778 3110
rect 6436 2272 7084 6802
rect 9172 6774 11542 6784
rect 9172 6672 11540 6682
rect 9172 6592 11540 6602
rect 9172 6492 11542 6502
rect 9172 6418 11542 6428
rect 9172 6316 11540 6326
rect 9172 6236 11540 6246
rect 9172 6136 11542 6146
rect 9172 6062 11542 6072
rect 9170 5960 11538 5970
rect 9170 5880 11538 5890
rect 9172 5778 11542 5788
rect 9172 5704 11542 5714
rect 9172 5604 11540 5614
rect 9172 5524 11540 5534
rect 9172 5422 11542 5432
rect 9172 5348 11542 5358
rect 9172 5246 11540 5256
rect 9172 5166 11540 5176
rect 9172 5066 11542 5076
rect 9172 4992 11542 5002
rect 9174 4892 11542 4902
rect 9172 4822 9174 4892
rect 9174 4812 11542 4822
rect 9172 4712 11542 4722
rect 9172 4638 11542 4648
rect 9172 4536 11540 4546
rect 9172 4456 11540 4466
rect 9172 4356 11542 4366
rect 9172 4282 11542 4292
rect 9172 4180 11540 4190
rect 9172 4100 11540 4110
rect 9172 3998 11542 4008
rect 9172 3924 11542 3934
rect 9172 3824 11540 3834
rect 9172 3744 11540 3754
rect 9172 3642 11542 3652
rect 9172 3568 11542 3578
rect 9172 3468 11540 3478
rect 9172 3388 11540 3398
rect 9172 3288 11542 3298
rect 9172 3214 11542 3224
rect 9172 3112 11540 3122
rect 9172 3032 11540 3042
rect 9172 2932 11542 2942
rect 9172 2858 11542 2868
rect 11594 2286 11754 20760
rect 11808 20730 14178 20740
rect 11808 20656 14178 20666
rect 14536 20728 16910 20738
rect 14536 20660 16910 20670
rect 11808 20556 14176 20566
rect 11808 20476 14176 20486
rect 14540 20558 16908 20568
rect 14540 20478 16908 20488
rect 11808 20374 14178 20384
rect 11808 20300 14178 20310
rect 14536 20372 16910 20382
rect 14536 20304 16910 20314
rect 11808 20200 14176 20210
rect 11808 20120 14176 20130
rect 14540 20200 16908 20210
rect 14540 20120 16908 20130
rect 11808 20018 14178 20028
rect 11808 19944 14178 19954
rect 14536 20016 16910 20026
rect 14536 19948 16910 19958
rect 11808 19844 14176 19854
rect 11808 19764 14176 19774
rect 14540 19844 16908 19854
rect 14540 19764 16908 19774
rect 11808 19662 14178 19672
rect 11808 19588 14178 19598
rect 14536 19660 16910 19670
rect 14536 19592 16910 19602
rect 11808 19488 14176 19498
rect 11808 19408 14176 19418
rect 14540 19486 16908 19496
rect 14540 19406 16908 19416
rect 11808 19308 14178 19318
rect 11808 19234 14178 19244
rect 14536 19304 16910 19314
rect 14536 19236 16910 19246
rect 11808 19132 14176 19142
rect 11808 19052 14176 19062
rect 14540 19132 16908 19142
rect 14540 19052 16908 19062
rect 11808 18950 14178 18960
rect 11808 18876 14178 18886
rect 14536 18948 16910 18958
rect 14536 18880 16910 18890
rect 11808 18776 14176 18786
rect 11808 18696 14176 18706
rect 14540 18776 16908 18786
rect 14540 18696 16908 18706
rect 11808 18594 14178 18604
rect 11808 18520 14178 18530
rect 14536 18592 16910 18602
rect 14536 18524 16910 18534
rect 11808 18420 14176 18430
rect 11808 18340 14176 18350
rect 14540 18420 16908 18430
rect 14540 18340 16908 18350
rect 11808 18238 14178 18248
rect 11808 18164 14178 18174
rect 14536 18236 16910 18246
rect 14536 18168 16910 18178
rect 11808 18064 14176 18074
rect 11808 17984 14176 17994
rect 14540 18064 16908 18074
rect 14540 17984 16908 17994
rect 11808 17882 14178 17892
rect 11808 17808 14178 17818
rect 14536 17880 16910 17890
rect 14536 17812 16910 17822
rect 11808 17708 14176 17718
rect 11808 17628 14176 17638
rect 14540 17708 16908 17718
rect 14540 17628 16908 17638
rect 11808 17528 14178 17538
rect 11808 17454 14178 17464
rect 14536 17524 16910 17534
rect 14536 17456 16910 17466
rect 11808 17352 14176 17362
rect 11808 17272 14176 17282
rect 14540 17352 16908 17362
rect 14540 17272 16908 17282
rect 11808 17172 14178 17182
rect 11808 17098 14178 17108
rect 14536 17168 16910 17178
rect 14536 17100 16910 17110
rect 11808 16996 14176 17006
rect 11808 16916 14176 16926
rect 14540 16996 16908 17006
rect 14540 16916 16908 16926
rect 11808 16816 14178 16826
rect 11808 16742 14178 16752
rect 14536 16812 16910 16822
rect 14536 16744 16910 16754
rect 11808 16640 14176 16650
rect 11808 16560 14176 16570
rect 14540 16640 16908 16650
rect 14540 16560 16908 16570
rect 11808 16460 14178 16470
rect 11808 16386 14178 16396
rect 14536 16456 16910 16466
rect 14536 16388 16910 16398
rect 11808 16286 14176 16296
rect 11808 16206 14176 16216
rect 14540 16284 16908 16294
rect 14540 16204 16908 16214
rect 11808 16102 14178 16112
rect 11808 16028 14178 16038
rect 14536 16100 16910 16110
rect 14536 16032 16910 16042
rect 11808 15928 14176 15938
rect 11808 15848 14176 15858
rect 14540 15926 16908 15936
rect 14540 15846 16908 15856
rect 11808 15746 14178 15756
rect 11808 15672 14178 15682
rect 14536 15744 16910 15754
rect 14536 15676 16910 15686
rect 11808 15572 14176 15582
rect 11808 15492 14176 15502
rect 14540 15572 16908 15582
rect 14540 15492 16908 15502
rect 11808 15392 14178 15402
rect 11808 15318 14178 15328
rect 14536 15388 16910 15398
rect 14536 15320 16910 15330
rect 11808 15216 14176 15226
rect 11808 15136 14176 15146
rect 14540 15216 16908 15226
rect 14540 15136 16908 15146
rect 11808 15034 14178 15044
rect 11808 14960 14178 14970
rect 14536 15032 16910 15042
rect 14536 14964 16910 14974
rect 11808 14860 14176 14870
rect 11808 14780 14176 14790
rect 14540 14860 16908 14870
rect 14540 14780 16908 14790
rect 11808 14680 14178 14690
rect 11808 14606 14178 14616
rect 14536 14676 16910 14686
rect 14536 14608 16910 14618
rect 11808 14504 14176 14514
rect 11808 14424 14176 14434
rect 14540 14504 16908 14514
rect 14540 14424 16908 14434
rect 11808 14322 14178 14332
rect 11808 14248 14178 14258
rect 14536 14320 16910 14330
rect 14536 14252 16910 14262
rect 11808 14148 14176 14158
rect 11808 14068 14176 14078
rect 14540 14146 16908 14156
rect 14540 14066 16908 14076
rect 11808 13968 14178 13978
rect 11808 13894 14178 13904
rect 14536 13964 16910 13974
rect 14536 13896 16910 13906
rect 11808 13792 14176 13802
rect 11808 13712 14176 13722
rect 14540 13792 16908 13802
rect 14540 13712 16908 13722
rect 11808 13612 14178 13622
rect 11808 13538 14178 13548
rect 14536 13608 16910 13618
rect 14536 13540 16910 13550
rect 11808 13436 14176 13446
rect 11808 13356 14176 13366
rect 14540 13436 16908 13446
rect 14540 13356 16908 13366
rect 11808 13254 14178 13264
rect 11808 13180 14178 13190
rect 14536 13252 16910 13262
rect 14536 13184 16910 13194
rect 11808 13080 14176 13090
rect 11808 13000 14176 13010
rect 14540 13080 16908 13090
rect 14540 13000 16908 13010
rect 11808 12898 14178 12908
rect 11808 12824 14178 12834
rect 14536 12896 16910 12906
rect 14536 12828 16910 12838
rect 11808 12724 14176 12734
rect 11808 12644 14176 12654
rect 14540 12724 16908 12734
rect 14540 12644 16908 12654
rect 11808 12544 14178 12554
rect 11808 12470 14178 12480
rect 14536 12540 16910 12550
rect 14536 12472 16910 12482
rect 11808 12368 14176 12378
rect 11808 12288 14176 12298
rect 14540 12368 16908 12378
rect 14540 12288 16908 12298
rect 11808 12186 14178 12196
rect 11808 12112 14178 12122
rect 14536 12184 16910 12194
rect 14536 12116 16910 12126
rect 11808 12012 14176 12022
rect 11808 11932 14176 11942
rect 14540 12012 16908 12022
rect 14540 11932 16908 11942
rect 11808 11830 14178 11840
rect 11808 11756 14178 11766
rect 14536 11828 16910 11838
rect 14536 11760 16910 11770
rect 11808 11656 14176 11666
rect 11808 11576 14176 11586
rect 14540 11656 16908 11666
rect 14540 11576 16908 11586
rect 11808 11476 14178 11486
rect 11808 11402 14178 11412
rect 14536 11472 16910 11482
rect 14536 11404 16910 11414
rect 11808 11300 14176 11310
rect 11808 11220 14176 11230
rect 14540 11300 16908 11310
rect 14540 11220 16908 11230
rect 11808 11120 14178 11130
rect 11808 11046 14178 11056
rect 14536 11116 16910 11126
rect 14536 11048 16910 11058
rect 11808 10944 14176 10954
rect 11808 10864 14176 10874
rect 14540 10946 16908 10956
rect 14540 10866 16908 10876
rect 11808 10764 14178 10774
rect 11808 10690 14178 10700
rect 14536 10760 16910 10770
rect 14536 10692 16910 10702
rect 11808 10588 14176 10598
rect 11808 10508 14176 10518
rect 14538 10586 16906 10596
rect 14538 10506 16906 10516
rect 11808 10408 14178 10418
rect 11808 10334 14178 10344
rect 14536 10404 16910 10414
rect 14536 10336 16910 10346
rect 11808 10232 14176 10242
rect 11808 10152 14176 10162
rect 14540 10232 16908 10242
rect 14540 10152 16908 10162
rect 11808 10052 14178 10062
rect 11808 9978 14178 9988
rect 14536 10048 16910 10058
rect 14536 9980 16910 9990
rect 11808 9876 14176 9886
rect 11808 9796 14176 9806
rect 14540 9876 16908 9886
rect 14540 9796 16908 9806
rect 11808 9696 14178 9706
rect 11808 9622 14178 9632
rect 14536 9692 16910 9702
rect 14536 9624 16910 9634
rect 11808 9520 14176 9530
rect 11808 9440 14176 9450
rect 14538 9520 16906 9530
rect 14538 9440 16906 9450
rect 11808 9340 14178 9350
rect 11808 9266 14178 9276
rect 14536 9338 16910 9348
rect 14536 9270 16910 9280
rect 11810 9164 14178 9174
rect 11810 9084 14178 9094
rect 14538 9164 16906 9174
rect 14538 9084 16906 9094
rect 11808 8982 14178 8992
rect 11808 8908 14178 8918
rect 14536 8980 16910 8990
rect 14536 8912 16910 8922
rect 11810 8808 14178 8818
rect 11810 8728 14178 8738
rect 14538 8806 16906 8816
rect 14538 8726 16906 8736
rect 11808 8628 14178 8638
rect 11808 8554 14178 8564
rect 14534 8624 16908 8634
rect 14534 8556 16908 8566
rect 11808 8452 14176 8462
rect 11808 8372 14176 8382
rect 14538 8452 16906 8462
rect 14538 8372 16906 8382
rect 11806 8272 14176 8282
rect 11806 8198 14176 8208
rect 14536 8268 16910 8278
rect 14536 8200 16910 8210
rect 11810 8096 14178 8106
rect 11810 8016 14178 8026
rect 14540 8096 16908 8106
rect 14540 8016 16908 8026
rect 11808 7914 14178 7924
rect 11808 7840 14178 7850
rect 14536 7912 16910 7922
rect 14536 7844 16910 7854
rect 11808 7740 14176 7750
rect 11808 7660 14176 7670
rect 14540 7742 16908 7752
rect 14540 7662 16908 7672
rect 11808 7560 14178 7570
rect 11808 7486 14178 7496
rect 14536 7556 16910 7566
rect 14536 7488 16910 7498
rect 11808 7384 14176 7394
rect 11808 7304 14176 7314
rect 14540 7384 16908 7394
rect 14540 7304 16908 7314
rect 11808 7204 14178 7214
rect 11808 7130 14178 7140
rect 14536 7200 16910 7210
rect 14536 7132 16910 7142
rect 11810 7028 14178 7038
rect 11810 6948 14178 6958
rect 14540 7026 16908 7036
rect 14540 6946 16908 6956
rect 11808 6848 14178 6858
rect 11808 6774 14178 6784
rect 14536 6844 16910 6854
rect 14536 6776 16910 6786
rect 11808 6672 14176 6682
rect 11808 6592 14176 6602
rect 14540 6672 16908 6682
rect 14540 6592 16908 6602
rect 11808 6490 14178 6500
rect 11808 6416 14178 6426
rect 14536 6488 16910 6498
rect 14536 6420 16910 6430
rect 11810 6316 14178 6326
rect 11810 6236 14178 6246
rect 14540 6316 16908 6326
rect 14540 6236 16908 6246
rect 11808 6136 14178 6146
rect 11808 6062 14178 6072
rect 14536 6132 16910 6142
rect 14536 6064 16910 6074
rect 11810 5960 14178 5970
rect 11810 5880 14178 5890
rect 14540 5962 16908 5972
rect 14540 5882 16908 5892
rect 11808 5778 14178 5788
rect 11808 5704 14178 5714
rect 14536 5776 16910 5786
rect 14536 5708 16910 5718
rect 11808 5604 14176 5614
rect 11808 5524 14176 5534
rect 14540 5604 16908 5614
rect 14540 5524 16908 5534
rect 11808 5422 14178 5432
rect 11808 5348 14178 5358
rect 14536 5420 16910 5430
rect 14536 5352 16910 5362
rect 11808 5248 14176 5258
rect 11808 5168 14176 5178
rect 14540 5246 16908 5256
rect 14540 5166 16908 5176
rect 11806 5066 14176 5076
rect 11806 4992 14176 5002
rect 14536 5064 16910 5074
rect 14536 4996 16910 5006
rect 11808 4892 14176 4902
rect 11808 4812 14176 4822
rect 14540 4892 16908 4902
rect 14540 4812 16908 4822
rect 11806 4712 14176 4722
rect 11806 4638 14176 4648
rect 14536 4708 16910 4718
rect 14536 4640 16910 4650
rect 11808 4536 14176 4546
rect 11808 4456 14176 4466
rect 14540 4536 16908 4546
rect 14540 4456 16908 4466
rect 11808 4354 14178 4364
rect 11808 4280 14178 4290
rect 14536 4352 16910 4362
rect 14536 4284 16910 4294
rect 11808 4180 14176 4190
rect 11808 4100 14176 4110
rect 14540 4180 16908 4190
rect 14540 4100 16908 4110
rect 11808 3998 14178 4008
rect 11808 3924 14178 3934
rect 14536 3996 16910 4006
rect 14536 3928 16910 3938
rect 11808 3824 14176 3834
rect 11808 3744 14176 3754
rect 14540 3824 16908 3834
rect 14540 3744 16908 3754
rect 11806 3642 14176 3652
rect 11806 3568 14176 3578
rect 14536 3640 16910 3650
rect 14536 3572 16910 3582
rect 11808 3468 14176 3478
rect 11808 3388 14176 3398
rect 14540 3466 16908 3476
rect 14540 3386 16908 3396
rect 11808 3288 14178 3298
rect 11808 3214 14178 3224
rect 14536 3284 16910 3294
rect 14536 3216 16910 3226
rect 11808 3112 14176 3122
rect 11808 3032 14176 3042
rect 14540 3112 16908 3122
rect 14540 3032 16908 3042
rect 11806 2932 14176 2942
rect 11806 2858 14176 2868
rect 14536 2928 16910 2938
rect 14536 2860 16910 2870
rect 16962 2286 17122 20760
rect 17172 20728 19546 20738
rect 17172 20660 19546 20670
rect 17176 20556 19544 20566
rect 17176 20476 19544 20486
rect 17172 20372 19546 20382
rect 17172 20304 19546 20314
rect 17176 20200 19544 20210
rect 17176 20120 19544 20130
rect 17172 20016 19546 20026
rect 17172 19948 19546 19958
rect 17176 19844 19544 19854
rect 17176 19764 19544 19774
rect 17172 19660 19546 19670
rect 17172 19592 19546 19602
rect 17176 19486 19544 19496
rect 17176 19406 19544 19416
rect 17172 19304 19546 19314
rect 17172 19236 19546 19246
rect 17176 19132 19544 19142
rect 17176 19052 19544 19062
rect 17172 18948 19546 18958
rect 17172 18880 19546 18890
rect 17176 18776 19544 18786
rect 17176 18696 19544 18706
rect 17172 18592 19546 18602
rect 17172 18524 19546 18534
rect 17176 18420 19544 18430
rect 17176 18340 19544 18350
rect 17172 18236 19546 18246
rect 17172 18168 19546 18178
rect 17176 18064 19544 18074
rect 17176 17984 19544 17994
rect 17172 17880 19546 17890
rect 17172 17812 19546 17822
rect 17176 17706 19544 17716
rect 17176 17626 19544 17636
rect 17172 17524 19546 17534
rect 17172 17456 19546 17466
rect 17176 17352 19544 17362
rect 17176 17272 19544 17282
rect 17172 17168 19546 17178
rect 17172 17100 19546 17110
rect 17176 16996 19544 17006
rect 17176 16916 19544 16926
rect 17172 16812 19546 16822
rect 17172 16744 19546 16754
rect 17176 16640 19544 16650
rect 17176 16560 19544 16570
rect 17172 16456 19546 16466
rect 17172 16388 19546 16398
rect 17176 16284 19544 16294
rect 17176 16204 19544 16214
rect 17172 16100 19546 16110
rect 17172 16032 19546 16042
rect 17176 15928 19544 15938
rect 17176 15848 19544 15858
rect 17172 15744 19546 15754
rect 17172 15676 19546 15686
rect 17176 15572 19544 15582
rect 17176 15492 19544 15502
rect 17172 15388 19546 15398
rect 17172 15320 19546 15330
rect 17176 15216 19544 15226
rect 17176 15136 19544 15146
rect 17172 15032 19546 15042
rect 17172 14964 19546 14974
rect 17176 14860 19544 14870
rect 17176 14780 19544 14790
rect 17172 14676 19546 14686
rect 17172 14608 19546 14618
rect 17176 14504 19544 14514
rect 17176 14424 19544 14434
rect 17172 14318 19546 14328
rect 17172 14250 19546 14260
rect 20904 14194 20926 25168
rect 21000 14194 21010 25168
rect 21052 25160 23024 25170
rect 21054 25056 23024 25066
rect 21054 24982 23024 24992
rect 21052 24872 23024 24882
rect 21052 24806 23024 24816
rect 21054 24700 23024 24710
rect 21054 24626 23024 24636
rect 21052 24516 23024 24526
rect 21052 24450 23024 24460
rect 21054 24342 23024 24352
rect 21054 24268 23024 24278
rect 21052 24160 23024 24170
rect 21052 24094 23024 24104
rect 21054 23986 23024 23996
rect 21054 23912 23024 23922
rect 21052 23804 23024 23814
rect 21052 23738 23024 23748
rect 21052 23632 23022 23642
rect 21052 23558 23022 23568
rect 21052 23448 23024 23458
rect 21052 23382 23024 23392
rect 21054 23274 23024 23284
rect 21054 23200 23024 23210
rect 21052 23092 23024 23102
rect 21052 23026 23024 23036
rect 21054 22920 23024 22930
rect 21054 22846 23024 22856
rect 21052 22736 23024 22746
rect 21052 22670 23024 22680
rect 21054 22562 23024 22572
rect 21054 22488 23024 22498
rect 21052 22380 23024 22390
rect 21052 22314 23024 22324
rect 21054 22206 23024 22216
rect 21054 22132 23024 22142
rect 21052 22024 23024 22034
rect 21052 21958 23024 21968
rect 21054 21852 23024 21862
rect 21054 21778 23024 21788
rect 21052 21668 23024 21678
rect 21052 21602 23024 21612
rect 21054 21494 23024 21504
rect 21054 21420 23024 21430
rect 21052 21312 23024 21322
rect 21052 21246 23024 21256
rect 21054 21140 23024 21150
rect 21054 21066 23024 21076
rect 21052 20956 23024 20966
rect 21052 20890 23024 20900
rect 21052 20782 23022 20792
rect 21052 20708 23022 20718
rect 21052 20600 23024 20610
rect 21052 20534 23024 20544
rect 21054 20424 23024 20434
rect 21054 20350 23024 20360
rect 21052 20244 23024 20254
rect 21052 20178 23024 20188
rect 21052 20072 23022 20082
rect 21052 19998 23022 20008
rect 21052 19888 23024 19898
rect 21052 19822 23024 19832
rect 21054 19714 23024 19724
rect 21054 19640 23024 19650
rect 21052 19532 23024 19542
rect 21052 19466 23024 19476
rect 21052 19360 23022 19370
rect 21052 19286 23022 19296
rect 21052 19176 23024 19186
rect 21052 19110 23024 19120
rect 21054 19002 23024 19012
rect 21054 18928 23024 18938
rect 21052 18820 23024 18830
rect 21052 18754 23024 18764
rect 21052 18646 23022 18656
rect 21052 18572 23022 18582
rect 21052 18464 23024 18474
rect 21052 18398 23024 18408
rect 21054 18290 23024 18300
rect 21054 18216 23024 18226
rect 21052 18108 23024 18118
rect 21052 18042 23024 18052
rect 21054 17934 23024 17944
rect 21054 17860 23024 17870
rect 21052 17752 23024 17762
rect 21052 17686 23024 17696
rect 21054 17578 23024 17588
rect 21054 17504 23024 17514
rect 21052 17396 23024 17406
rect 21052 17330 23024 17340
rect 21054 17222 23024 17232
rect 21054 17148 23024 17158
rect 21052 17040 23024 17050
rect 21052 16974 23024 16984
rect 21054 16866 23024 16876
rect 21054 16792 23024 16802
rect 21052 16684 23024 16694
rect 21052 16618 23024 16628
rect 21052 16510 23022 16520
rect 21052 16436 23022 16446
rect 21052 16328 23024 16338
rect 21052 16262 23024 16272
rect 21054 16154 23024 16164
rect 21054 16080 23024 16090
rect 21052 15972 23024 15982
rect 21052 15906 23024 15916
rect 21054 15800 23024 15810
rect 21054 15726 23024 15736
rect 21052 15616 23024 15626
rect 21052 15550 23024 15560
rect 21054 15442 23024 15452
rect 21054 15368 23024 15378
rect 21052 15260 23024 15270
rect 21052 15194 23024 15204
rect 21054 15086 23024 15096
rect 21054 15012 23024 15022
rect 21052 14904 23024 14914
rect 21052 14838 23024 14848
rect 21054 14732 23024 14742
rect 21054 14658 23024 14668
rect 21052 14548 23024 14558
rect 21052 14482 23024 14492
rect 21054 14374 23024 14384
rect 21054 14300 23024 14310
rect 17176 14148 19544 14158
rect 20904 14132 21006 14194
rect 21052 14192 23024 14202
rect 21052 14126 23024 14136
rect 17176 14068 19544 14078
rect 17172 13964 19546 13974
rect 17172 13896 19546 13906
rect 21052 13968 23024 13978
rect 21052 13900 23024 13910
rect 17176 13792 19544 13802
rect 17176 13712 19544 13722
rect 21052 13788 23024 13798
rect 21052 13720 23024 13730
rect 17172 13608 19546 13618
rect 17172 13540 19546 13550
rect 21052 13610 23024 13620
rect 21052 13542 23024 13552
rect 17176 13436 19544 13446
rect 17176 13356 19544 13366
rect 21052 13432 23024 13442
rect 21052 13364 23024 13374
rect 17172 13252 19546 13262
rect 17172 13184 19546 13194
rect 21052 13254 23024 13264
rect 21052 13186 23024 13196
rect 17176 13080 19544 13090
rect 17176 13000 19544 13010
rect 21052 13076 23024 13086
rect 21052 13008 23024 13018
rect 17172 12896 19546 12906
rect 17172 12828 19546 12838
rect 21052 12898 23024 12908
rect 21052 12830 23024 12840
rect 17176 12724 19544 12734
rect 17176 12644 19544 12654
rect 21052 12720 23024 12730
rect 21052 12652 23024 12662
rect 17172 12540 19546 12550
rect 17172 12472 19546 12482
rect 21052 12542 23024 12552
rect 21052 12474 23024 12484
rect 17178 12368 19546 12378
rect 17178 12288 19546 12298
rect 21052 12364 23024 12374
rect 21052 12296 23024 12306
rect 17172 12184 19546 12194
rect 17172 12116 19546 12126
rect 21052 12186 23024 12196
rect 21052 12118 23024 12128
rect 17178 12012 19546 12022
rect 17178 11932 19546 11942
rect 21052 12008 23024 12018
rect 21052 11940 23024 11950
rect 17172 11828 19546 11838
rect 17172 11760 19546 11770
rect 21052 11830 23024 11840
rect 21052 11762 23024 11772
rect 17176 11656 19544 11666
rect 17176 11576 19544 11586
rect 21052 11652 23024 11662
rect 21052 11584 23024 11594
rect 17172 11472 19546 11482
rect 17172 11404 19546 11414
rect 21052 11474 23024 11484
rect 21052 11406 23024 11416
rect 17176 11300 19544 11310
rect 17176 11220 19544 11230
rect 21052 11296 23024 11306
rect 21052 11228 23024 11238
rect 17172 11116 19546 11126
rect 17172 11048 19546 11058
rect 21052 11118 23024 11128
rect 21052 11050 23024 11060
rect 17176 10944 19544 10954
rect 17176 10864 19544 10874
rect 21052 10940 23024 10950
rect 21052 10872 23024 10882
rect 17172 10760 19546 10770
rect 17172 10692 19546 10702
rect 21052 10762 23024 10772
rect 21052 10694 23024 10704
rect 17176 10588 19544 10598
rect 17176 10508 19544 10518
rect 21052 10584 23024 10594
rect 21052 10516 23024 10526
rect 17172 10404 19546 10414
rect 17172 10336 19546 10346
rect 21052 10406 23024 10416
rect 21052 10338 23024 10348
rect 17176 10232 19544 10242
rect 17176 10152 19544 10162
rect 21052 10228 23024 10238
rect 21052 10160 23024 10170
rect 17172 10048 19546 10058
rect 17172 9980 19546 9990
rect 21052 10050 23024 10060
rect 21052 9982 23024 9992
rect 17176 9876 19544 9886
rect 17176 9796 19544 9806
rect 21052 9872 23024 9882
rect 21052 9804 23024 9814
rect 17172 9692 19546 9702
rect 17172 9624 19546 9634
rect 21052 9694 23024 9704
rect 21052 9626 23024 9636
rect 17176 9520 19544 9530
rect 17176 9440 19544 9450
rect 21052 9516 23024 9526
rect 21052 9448 23024 9458
rect 17172 9336 19546 9346
rect 17172 9268 19546 9278
rect 21052 9338 23024 9348
rect 21052 9270 23024 9280
rect 17176 9164 19544 9174
rect 17176 9084 19544 9094
rect 21052 9160 23024 9170
rect 21052 9092 23024 9102
rect 17172 8980 19546 8990
rect 17172 8912 19546 8922
rect 21052 8982 23024 8992
rect 21052 8914 23024 8924
rect 17176 8808 19544 8818
rect 17176 8728 19544 8738
rect 21052 8804 23024 8814
rect 21052 8736 23024 8746
rect 17172 8624 19546 8634
rect 17172 8556 19546 8566
rect 21052 8626 23024 8636
rect 21052 8558 23024 8568
rect 17176 8452 19544 8462
rect 17176 8372 19544 8382
rect 21054 8448 23026 8458
rect 21054 8380 23026 8390
rect 17172 8268 19546 8278
rect 17172 8200 19546 8210
rect 21052 8270 23024 8280
rect 21052 8202 23024 8212
rect 17176 8096 19544 8106
rect 17176 8016 19544 8026
rect 21052 8092 23024 8102
rect 21052 8024 23024 8034
rect 17172 7912 19546 7922
rect 17172 7844 19546 7854
rect 21052 7914 23024 7924
rect 21052 7846 23024 7856
rect 17176 7740 19544 7750
rect 17176 7660 19544 7670
rect 21052 7736 23024 7746
rect 21052 7668 23024 7678
rect 17172 7556 19546 7566
rect 17172 7488 19546 7498
rect 21052 7558 23024 7568
rect 21052 7490 23024 7500
rect 17176 7384 19544 7394
rect 17176 7304 19544 7314
rect 21052 7380 23024 7390
rect 21052 7312 23024 7322
rect 17172 7198 19546 7208
rect 17172 7130 19546 7140
rect 21052 7202 23024 7212
rect 21052 7134 23024 7144
rect 17176 7028 19544 7038
rect 17176 6948 19544 6958
rect 21052 7024 23024 7034
rect 21052 6956 23024 6966
rect 17172 6844 19546 6854
rect 17172 6776 19546 6786
rect 21052 6848 23024 6858
rect 21052 6780 23024 6790
rect 17176 6672 19544 6682
rect 17176 6592 19544 6602
rect 21052 6668 23024 6678
rect 21052 6600 23024 6610
rect 17172 6488 19546 6498
rect 17172 6420 19546 6430
rect 21052 6490 23024 6500
rect 21052 6422 23024 6432
rect 17176 6316 19544 6326
rect 17176 6236 19544 6246
rect 21052 6312 23024 6322
rect 21052 6244 23024 6254
rect 17172 6132 19546 6142
rect 17172 6064 19546 6074
rect 21052 6134 23024 6144
rect 21052 6066 23024 6076
rect 17176 5960 19544 5970
rect 17176 5880 19544 5890
rect 21052 5956 23024 5966
rect 21052 5888 23024 5898
rect 17172 5776 19546 5786
rect 17172 5708 19546 5718
rect 21052 5778 23024 5788
rect 21052 5710 23024 5720
rect 17176 5604 19544 5614
rect 17176 5524 19544 5534
rect 21052 5600 23024 5610
rect 21052 5532 23024 5542
rect 17172 5420 19546 5430
rect 17172 5352 19546 5362
rect 21052 5422 23024 5432
rect 21052 5354 23024 5364
rect 17176 5248 19544 5258
rect 17176 5168 19544 5178
rect 21052 5244 23024 5254
rect 21052 5176 23024 5186
rect 17172 5064 19546 5074
rect 17172 4996 19546 5006
rect 21052 5068 23024 5078
rect 21052 5000 23024 5010
rect 17176 4892 19544 4902
rect 17176 4812 19544 4822
rect 21052 4888 23024 4898
rect 21052 4820 23024 4830
rect 17172 4708 19546 4718
rect 17172 4640 19546 4650
rect 21052 4710 23024 4720
rect 21052 4642 23024 4652
rect 17176 4536 19544 4546
rect 17176 4456 19544 4466
rect 21052 4532 23024 4542
rect 21052 4464 23024 4474
rect 17172 4352 19546 4362
rect 17172 4284 19546 4294
rect 21052 4354 23024 4364
rect 21052 4286 23024 4296
rect 17176 4180 19544 4190
rect 17176 4100 19544 4110
rect 21052 4176 23024 4186
rect 21052 4108 23024 4118
rect 17172 3994 19546 4004
rect 17172 3926 19546 3936
rect 21052 4000 23024 4010
rect 21052 3932 23024 3942
rect 17176 3824 19544 3834
rect 17176 3744 19544 3754
rect 21052 3820 23024 3830
rect 21052 3752 23024 3762
rect 17172 3640 19546 3650
rect 17172 3572 19546 3582
rect 21052 3642 23024 3652
rect 21052 3574 23024 3584
rect 17176 3468 19544 3478
rect 17176 3388 19544 3398
rect 21052 3464 23024 3474
rect 21052 3396 23024 3406
rect 17170 3284 19544 3294
rect 17170 3216 19544 3226
rect 21052 3286 23024 3296
rect 21052 3218 23024 3228
rect 17176 3112 19544 3122
rect 17176 3032 19544 3042
rect 21052 3108 23024 3118
rect 21052 3040 23024 3050
rect 17170 2928 19544 2938
rect 17170 2860 19544 2870
rect 21052 2930 23024 2940
rect 21052 2862 23024 2872
rect 23068 2840 23170 25240
rect 25106 2734 25116 40588
rect 25640 2734 25650 40588
rect 25110 2722 25646 2734
rect 6232 1280 6242 2272
rect 7252 1280 7262 2272
rect 11172 1294 11182 2286
rect 12192 1294 12202 2286
rect 16514 1294 16524 2286
rect 17534 1294 17544 2286
<< via1 >>
rect 23738 43240 27086 43860
rect 3018 38138 4792 38204
rect 3012 38026 4800 38080
rect 3018 37902 4792 37968
rect 3012 37790 4800 37844
rect 3018 37666 4792 37732
rect 3012 37554 4800 37608
rect 3018 37430 4792 37496
rect 3012 37318 4800 37372
rect 3018 37194 4792 37260
rect 3012 37082 4800 37136
rect 3018 36958 4792 37024
rect 3012 36846 4800 36900
rect 3018 36722 4792 36788
rect 3012 36610 4800 36664
rect 3018 36486 4792 36552
rect 3012 36374 4800 36428
rect 3018 36250 4792 36316
rect 3012 36138 4800 36192
rect 3018 36014 4792 36080
rect 3012 35902 4800 35956
rect 3018 35778 4792 35844
rect 3012 35666 4800 35720
rect 3018 35542 4792 35608
rect 3012 35430 4800 35484
rect 3018 35306 4792 35372
rect 3012 35194 4800 35248
rect 3018 35070 4792 35136
rect 3012 34958 4800 35012
rect 3018 34834 4792 34900
rect 3012 34722 4800 34776
rect 3018 34598 4792 34664
rect 3012 34486 4800 34540
rect 3018 34362 4792 34428
rect 3012 34250 4800 34304
rect 3018 34126 4792 34192
rect 3012 34014 4800 34068
rect 3018 33890 4792 33956
rect 3012 33778 4800 33832
rect 3018 33654 4792 33720
rect 3012 33542 4800 33596
rect 3018 33418 4792 33484
rect 3012 33306 4800 33360
rect 3018 33182 4792 33248
rect 3012 33070 4800 33124
rect 3018 32946 4792 33012
rect 3012 32834 4800 32888
rect 3018 32710 4792 32776
rect 3012 32598 4800 32652
rect 3018 32474 4792 32540
rect 3012 32362 4800 32416
rect 3018 32238 4792 32304
rect 3012 32126 4800 32180
rect 3018 32002 4792 32068
rect 3012 31890 4800 31944
rect 3016 31766 4790 31832
rect 3012 31654 4800 31708
rect 3018 31530 4792 31596
rect 3012 31418 4800 31472
rect 3018 31294 4792 31360
rect 3012 31182 4800 31236
rect 3018 31060 4792 31120
rect 2784 3110 3772 29890
rect 20656 40396 23026 40460
rect 20658 40280 23028 40338
rect 20656 40160 23026 40224
rect 20656 40046 23026 40104
rect 20654 39924 23024 39988
rect 20658 39806 23028 39864
rect 20654 39688 23024 39752
rect 20656 39574 23026 39632
rect 20656 39452 23026 39516
rect 20656 39336 23026 39394
rect 20654 39214 23024 39278
rect 20656 39102 23026 39160
rect 20656 38978 23026 39042
rect 20656 38866 23026 38924
rect 20654 38746 23024 38810
rect 20658 38628 23028 38686
rect 20656 38506 23026 38570
rect 20656 38392 23026 38450
rect 20654 38270 23024 38334
rect 20656 38156 23026 38214
rect 20654 38034 23024 38098
rect 20656 37920 23026 37978
rect 20656 37798 23026 37862
rect 20658 37686 23028 37744
rect 20656 37562 23026 37626
rect 20656 37448 23026 37506
rect 20656 37326 23026 37390
rect 20658 37210 23028 37268
rect 20654 37092 23024 37156
rect 20658 36976 23028 37034
rect 20658 36856 23028 36920
rect 20658 36740 23028 36798
rect 20656 36618 23026 36682
rect 20656 36504 23026 36562
rect 20658 36382 23028 36446
rect 20658 36268 23028 36326
rect 20658 36146 23028 36210
rect 20656 36032 23026 36090
rect 20658 35912 23028 35976
rect 20656 35798 23026 35856
rect 20654 35674 23024 35738
rect 20658 35562 23028 35620
rect 20654 35436 23024 35500
rect 20656 35326 23026 35384
rect 20656 35202 23026 35266
rect 20656 35090 23026 35148
rect 20656 34966 23026 35030
rect 20656 34852 23026 34910
rect 20658 34730 23028 34794
rect 20658 34616 23028 34674
rect 20654 34496 23024 34560
rect 20660 34380 23030 34438
rect 20654 34258 23024 34322
rect 20658 34144 23028 34202
rect 20656 34024 23026 34088
rect 20656 33906 23026 33964
rect 20656 33786 23026 33850
rect 20656 33674 23026 33732
rect 20656 33550 23026 33614
rect 20656 33436 23026 33494
rect 20656 33316 23026 33380
rect 20658 33202 23028 33260
rect 20656 33080 23026 33144
rect 20658 32964 23028 33022
rect 20656 32842 23026 32906
rect 20656 32730 23026 32788
rect 20658 32608 23028 32672
rect 20656 32494 23026 32552
rect 20658 32374 23028 32438
rect 20656 32256 23026 32314
rect 20656 32134 23026 32198
rect 20656 32020 23026 32078
rect 20656 31900 23026 31964
rect 20658 31782 23028 31840
rect 20656 31662 23026 31726
rect 20658 31548 23028 31606
rect 20656 31428 23026 31492
rect 20658 31314 23028 31372
rect 20656 31192 23026 31256
rect 20656 31076 23026 31134
rect 20654 30956 23024 31020
rect 20656 30842 23026 30900
rect 20656 30718 23026 30782
rect 20656 30604 23026 30662
rect 20656 30482 23026 30546
rect 20656 30368 23026 30426
rect 20656 30248 23026 30312
rect 20658 30130 23028 30188
rect 20656 30010 23026 30074
rect 20658 29896 23028 29954
rect 20658 29776 23028 29840
rect 18478 22294 18982 22684
rect 19814 22660 19974 22772
rect 21052 25170 23024 25226
rect 19810 21030 19970 21144
rect 9172 20666 11542 20730
rect 9174 20486 11542 20556
rect 9172 20310 11542 20374
rect 9172 20130 11540 20200
rect 9172 19954 11542 20018
rect 9172 19774 11540 19844
rect 9172 19598 11542 19662
rect 9172 19420 11540 19490
rect 9172 19244 11542 19308
rect 9172 19062 11540 19132
rect 9172 18886 11542 18950
rect 9172 18706 11540 18776
rect 9172 18530 11542 18594
rect 9172 18350 11540 18420
rect 9172 18174 11542 18238
rect 9172 17994 11540 18064
rect 9172 17818 11542 17882
rect 9172 17638 11540 17708
rect 9172 17464 11542 17528
rect 9172 17280 11540 17350
rect 9172 17108 11542 17172
rect 9172 16926 11540 16996
rect 9172 16752 11542 16816
rect 9172 16570 11540 16640
rect 9172 16398 11542 16462
rect 9172 16216 11540 16286
rect 9172 16038 11542 16102
rect 9172 15858 11540 15928
rect 4780 15648 6568 15710
rect 4782 15534 6570 15588
rect 4780 15412 6568 15474
rect 4782 15298 6570 15352
rect 4780 15176 6568 15238
rect 4782 15062 6570 15116
rect 4780 14940 6568 15002
rect 4782 14826 6570 14880
rect 4780 14704 6568 14766
rect 4782 14590 6570 14644
rect 4780 14468 6568 14530
rect 4782 14354 6570 14408
rect 4780 14232 6568 14294
rect 4780 14118 6568 14172
rect 4778 13996 6566 14058
rect 4780 13882 6568 13936
rect 4780 13760 6568 13822
rect 4782 13646 6570 13700
rect 4780 13524 6568 13586
rect 4782 13410 6570 13464
rect 4780 13288 6568 13350
rect 4782 13174 6570 13228
rect 4780 13052 6568 13114
rect 4782 12938 6570 12992
rect 4780 12816 6568 12878
rect 4782 12702 6570 12756
rect 4778 12580 6566 12642
rect 4782 12466 6570 12520
rect 4780 12344 6568 12406
rect 4782 12230 6570 12284
rect 4780 12108 6568 12170
rect 4782 11994 6570 12048
rect 4780 11872 6568 11934
rect 4782 11758 6570 11812
rect 4778 11636 6566 11698
rect 4782 11522 6570 11576
rect 4778 11400 6566 11462
rect 4782 11286 6570 11340
rect 4780 11164 6568 11226
rect 4782 11050 6570 11104
rect 4780 10928 6568 10990
rect 4782 10814 6570 10868
rect 4780 10692 6568 10754
rect 4782 10578 6570 10632
rect 4780 10456 6568 10518
rect 4782 10342 6570 10396
rect 4778 10220 6566 10282
rect 4782 10106 6570 10160
rect 4778 9984 6566 10046
rect 4782 9870 6570 9924
rect 4780 9748 6568 9810
rect 4782 9634 6570 9688
rect 4778 9512 6566 9574
rect 4782 9398 6570 9452
rect 4780 9276 6568 9338
rect 4780 9162 6568 9216
rect 4778 9038 6566 9100
rect 4780 8926 6568 8980
rect 4778 8804 6566 8866
rect 4780 8690 6568 8744
rect 4780 8568 6568 8630
rect 9172 15682 11542 15746
rect 9172 15502 11540 15572
rect 9172 15328 11542 15392
rect 9172 15146 11540 15216
rect 9172 14970 11542 15034
rect 9172 14790 11540 14860
rect 9172 14616 11542 14680
rect 9172 14434 11540 14504
rect 9172 14258 11542 14322
rect 9172 14078 11540 14148
rect 9172 13904 11542 13968
rect 9172 13722 11540 13792
rect 9172 13550 11542 13614
rect 9172 13366 11540 13436
rect 9172 13192 11542 13256
rect 9172 13010 11540 13080
rect 9172 12834 11542 12898
rect 9172 12654 11540 12724
rect 9172 12480 11542 12544
rect 9172 12298 11540 12368
rect 9172 12122 11542 12186
rect 9172 11942 11540 12012
rect 9172 11766 11542 11830
rect 9170 11586 11538 11656
rect 9172 11412 11542 11476
rect 9170 11230 11538 11300
rect 9172 11056 11542 11120
rect 9170 10874 11538 10944
rect 9172 10700 11542 10764
rect 9170 10518 11538 10588
rect 9170 10344 11540 10408
rect 9170 10160 11538 10230
rect 9172 9988 11542 10052
rect 9170 9806 11538 9876
rect 9172 9632 11542 9696
rect 9172 9450 11540 9520
rect 9172 9278 11542 9342
rect 9172 9094 11540 9164
rect 9172 8918 11542 8982
rect 9172 8736 11540 8806
rect 9172 8562 11542 8626
rect 9172 8382 11540 8452
rect 4788 8224 6568 8282
rect 9172 8208 11542 8272
rect 4788 7988 6568 8046
rect 9172 8026 11540 8096
rect 4788 7752 6568 7810
rect 9172 7852 11542 7916
rect 9172 7670 11540 7740
rect 9172 7496 11542 7560
rect 9172 7314 11540 7384
rect 9172 7140 11542 7204
rect 9172 6958 11540 7028
rect 9172 6784 11542 6848
rect 9172 6602 11540 6672
rect 9172 6428 11542 6492
rect 9172 6246 11540 6316
rect 9172 6072 11542 6136
rect 9170 5890 11538 5960
rect 9172 5714 11542 5778
rect 9172 5534 11540 5604
rect 9172 5358 11542 5422
rect 9172 5176 11540 5246
rect 9172 5002 11542 5066
rect 9174 4822 11542 4892
rect 9172 4648 11542 4712
rect 9172 4466 11540 4536
rect 9172 4292 11542 4356
rect 9172 4110 11540 4180
rect 9172 3934 11542 3998
rect 9172 3754 11540 3824
rect 9172 3578 11542 3642
rect 9172 3398 11540 3468
rect 9172 3224 11542 3288
rect 9172 3042 11540 3112
rect 9172 2868 11542 2932
rect 11808 20666 14178 20730
rect 14536 20670 16910 20728
rect 11808 20486 14176 20556
rect 14540 20488 16908 20558
rect 11808 20310 14178 20374
rect 14536 20314 16910 20372
rect 11808 20130 14176 20200
rect 14540 20130 16908 20200
rect 11808 19954 14178 20018
rect 14536 19958 16910 20016
rect 11808 19774 14176 19844
rect 14540 19774 16908 19844
rect 11808 19598 14178 19662
rect 14536 19602 16910 19660
rect 11808 19418 14176 19488
rect 14540 19416 16908 19486
rect 11808 19244 14178 19308
rect 14536 19246 16910 19304
rect 11808 19062 14176 19132
rect 14540 19062 16908 19132
rect 11808 18886 14178 18950
rect 14536 18890 16910 18948
rect 11808 18706 14176 18776
rect 14540 18706 16908 18776
rect 11808 18530 14178 18594
rect 14536 18534 16910 18592
rect 11808 18350 14176 18420
rect 14540 18350 16908 18420
rect 11808 18174 14178 18238
rect 14536 18178 16910 18236
rect 11808 17994 14176 18064
rect 14540 17994 16908 18064
rect 11808 17818 14178 17882
rect 14536 17822 16910 17880
rect 11808 17638 14176 17708
rect 14540 17638 16908 17708
rect 11808 17464 14178 17528
rect 14536 17466 16910 17524
rect 11808 17282 14176 17352
rect 14540 17282 16908 17352
rect 11808 17108 14178 17172
rect 14536 17110 16910 17168
rect 11808 16926 14176 16996
rect 14540 16926 16908 16996
rect 11808 16752 14178 16816
rect 14536 16754 16910 16812
rect 11808 16570 14176 16640
rect 14540 16570 16908 16640
rect 11808 16396 14178 16460
rect 14536 16398 16910 16456
rect 11808 16216 14176 16286
rect 14540 16214 16908 16284
rect 11808 16038 14178 16102
rect 14536 16042 16910 16100
rect 11808 15858 14176 15928
rect 14540 15856 16908 15926
rect 11808 15682 14178 15746
rect 14536 15686 16910 15744
rect 11808 15502 14176 15572
rect 14540 15502 16908 15572
rect 11808 15328 14178 15392
rect 14536 15330 16910 15388
rect 11808 15146 14176 15216
rect 14540 15146 16908 15216
rect 11808 14970 14178 15034
rect 14536 14974 16910 15032
rect 11808 14790 14176 14860
rect 14540 14790 16908 14860
rect 11808 14616 14178 14680
rect 14536 14618 16910 14676
rect 11808 14434 14176 14504
rect 14540 14434 16908 14504
rect 11808 14258 14178 14322
rect 14536 14262 16910 14320
rect 11808 14078 14176 14148
rect 14540 14076 16908 14146
rect 11808 13904 14178 13968
rect 14536 13906 16910 13964
rect 11808 13722 14176 13792
rect 14540 13722 16908 13792
rect 11808 13548 14178 13612
rect 14536 13550 16910 13608
rect 11808 13366 14176 13436
rect 14540 13366 16908 13436
rect 11808 13190 14178 13254
rect 14536 13194 16910 13252
rect 11808 13010 14176 13080
rect 14540 13010 16908 13080
rect 11808 12834 14178 12898
rect 14536 12838 16910 12896
rect 11808 12654 14176 12724
rect 14540 12654 16908 12724
rect 11808 12480 14178 12544
rect 14536 12482 16910 12540
rect 11808 12298 14176 12368
rect 14540 12298 16908 12368
rect 11808 12122 14178 12186
rect 14536 12126 16910 12184
rect 11808 11942 14176 12012
rect 14540 11942 16908 12012
rect 11808 11766 14178 11830
rect 14536 11770 16910 11828
rect 11808 11586 14176 11656
rect 14540 11586 16908 11656
rect 11808 11412 14178 11476
rect 14536 11414 16910 11472
rect 11808 11230 14176 11300
rect 14540 11230 16908 11300
rect 11808 11056 14178 11120
rect 14536 11058 16910 11116
rect 11808 10874 14176 10944
rect 14540 10876 16908 10946
rect 11808 10700 14178 10764
rect 14536 10702 16910 10760
rect 11808 10518 14176 10588
rect 14538 10516 16906 10586
rect 11808 10344 14178 10408
rect 14536 10346 16910 10404
rect 11808 10162 14176 10232
rect 14540 10162 16908 10232
rect 11808 9988 14178 10052
rect 14536 9990 16910 10048
rect 11808 9806 14176 9876
rect 14540 9806 16908 9876
rect 11808 9632 14178 9696
rect 14536 9634 16910 9692
rect 11808 9450 14176 9520
rect 14538 9450 16906 9520
rect 11808 9276 14178 9340
rect 14536 9280 16910 9338
rect 11810 9094 14178 9164
rect 14538 9094 16906 9164
rect 11808 8918 14178 8982
rect 14536 8922 16910 8980
rect 11810 8738 14178 8808
rect 14538 8736 16906 8806
rect 11808 8564 14178 8628
rect 14534 8566 16908 8624
rect 11808 8382 14176 8452
rect 14538 8382 16906 8452
rect 11806 8208 14176 8272
rect 14536 8210 16910 8268
rect 11810 8026 14178 8096
rect 14540 8026 16908 8096
rect 11808 7850 14178 7914
rect 14536 7854 16910 7912
rect 11808 7670 14176 7740
rect 14540 7672 16908 7742
rect 11808 7496 14178 7560
rect 14536 7498 16910 7556
rect 11808 7314 14176 7384
rect 14540 7314 16908 7384
rect 11808 7140 14178 7204
rect 14536 7142 16910 7200
rect 11810 6958 14178 7028
rect 14540 6956 16908 7026
rect 11808 6784 14178 6848
rect 14536 6786 16910 6844
rect 11808 6602 14176 6672
rect 14540 6602 16908 6672
rect 11808 6426 14178 6490
rect 14536 6430 16910 6488
rect 11810 6246 14178 6316
rect 14540 6246 16908 6316
rect 11808 6072 14178 6136
rect 14536 6074 16910 6132
rect 11810 5890 14178 5960
rect 14540 5892 16908 5962
rect 11808 5714 14178 5778
rect 14536 5718 16910 5776
rect 11808 5534 14176 5604
rect 14540 5534 16908 5604
rect 11808 5358 14178 5422
rect 14536 5362 16910 5420
rect 11808 5178 14176 5248
rect 14540 5176 16908 5246
rect 11806 5002 14176 5066
rect 14536 5006 16910 5064
rect 11808 4822 14176 4892
rect 14540 4822 16908 4892
rect 11806 4648 14176 4712
rect 14536 4650 16910 4708
rect 11808 4466 14176 4536
rect 14540 4466 16908 4536
rect 11808 4290 14178 4354
rect 14536 4294 16910 4352
rect 11808 4110 14176 4180
rect 14540 4110 16908 4180
rect 11808 3934 14178 3998
rect 14536 3938 16910 3996
rect 11808 3754 14176 3824
rect 14540 3754 16908 3824
rect 11806 3578 14176 3642
rect 14536 3582 16910 3640
rect 11808 3398 14176 3468
rect 14540 3396 16908 3466
rect 11808 3224 14178 3288
rect 14536 3226 16910 3284
rect 11808 3042 14176 3112
rect 14540 3042 16908 3112
rect 11806 2868 14176 2932
rect 14536 2870 16910 2928
rect 17172 20670 19546 20728
rect 17176 20486 19544 20556
rect 17172 20314 19546 20372
rect 17176 20130 19544 20200
rect 17172 19958 19546 20016
rect 17176 19774 19544 19844
rect 17172 19602 19546 19660
rect 17176 19416 19544 19486
rect 17172 19246 19546 19304
rect 17176 19062 19544 19132
rect 17172 18890 19546 18948
rect 17176 18706 19544 18776
rect 17172 18534 19546 18592
rect 17176 18350 19544 18420
rect 17172 18178 19546 18236
rect 17176 17994 19544 18064
rect 17172 17822 19546 17880
rect 17176 17636 19544 17706
rect 17172 17466 19546 17524
rect 17176 17282 19544 17352
rect 17172 17110 19546 17168
rect 17176 16926 19544 16996
rect 17172 16754 19546 16812
rect 17176 16570 19544 16640
rect 17172 16398 19546 16456
rect 17176 16214 19544 16284
rect 17172 16042 19546 16100
rect 17176 15858 19544 15928
rect 17172 15686 19546 15744
rect 17176 15502 19544 15572
rect 17172 15330 19546 15388
rect 17176 15146 19544 15216
rect 17172 14974 19546 15032
rect 17176 14790 19544 14860
rect 17172 14618 19546 14676
rect 17176 14434 19544 14504
rect 17172 14260 19546 14318
rect 20926 14194 21000 25168
rect 21054 24992 23024 25056
rect 21052 24816 23024 24872
rect 21054 24636 23024 24700
rect 21052 24460 23024 24516
rect 21054 24278 23024 24342
rect 21052 24104 23024 24160
rect 21054 23922 23024 23986
rect 21052 23748 23024 23804
rect 21052 23568 23022 23632
rect 21052 23392 23024 23448
rect 21054 23210 23024 23274
rect 21052 23036 23024 23092
rect 21054 22856 23024 22920
rect 21052 22680 23024 22736
rect 21054 22498 23024 22562
rect 21052 22324 23024 22380
rect 21054 22142 23024 22206
rect 21052 21968 23024 22024
rect 21054 21788 23024 21852
rect 21052 21612 23024 21668
rect 21054 21430 23024 21494
rect 21052 21256 23024 21312
rect 21054 21076 23024 21140
rect 21052 20900 23024 20956
rect 21052 20718 23022 20782
rect 21052 20544 23024 20600
rect 21054 20360 23024 20424
rect 21052 20188 23024 20244
rect 21052 20008 23022 20072
rect 21052 19832 23024 19888
rect 21054 19650 23024 19714
rect 21052 19476 23024 19532
rect 21052 19296 23022 19360
rect 21052 19120 23024 19176
rect 21054 18938 23024 19002
rect 21052 18764 23024 18820
rect 21052 18582 23022 18646
rect 21052 18408 23024 18464
rect 21054 18226 23024 18290
rect 21052 18052 23024 18108
rect 21054 17870 23024 17934
rect 21052 17696 23024 17752
rect 21054 17514 23024 17578
rect 21052 17340 23024 17396
rect 21054 17158 23024 17222
rect 21052 16984 23024 17040
rect 21054 16802 23024 16866
rect 21052 16628 23024 16684
rect 21052 16446 23022 16510
rect 21052 16272 23024 16328
rect 21054 16090 23024 16154
rect 21052 15916 23024 15972
rect 21054 15736 23024 15800
rect 21052 15560 23024 15616
rect 21054 15378 23024 15442
rect 21052 15204 23024 15260
rect 21054 15022 23024 15086
rect 21052 14848 23024 14904
rect 21054 14668 23024 14732
rect 21052 14492 23024 14548
rect 21054 14310 23024 14374
rect 17176 14078 19544 14148
rect 21052 14136 23024 14192
rect 17172 13906 19546 13964
rect 21052 13910 23024 13968
rect 17176 13722 19544 13792
rect 21052 13730 23024 13788
rect 17172 13550 19546 13608
rect 21052 13552 23024 13610
rect 17176 13366 19544 13436
rect 21052 13374 23024 13432
rect 17172 13194 19546 13252
rect 21052 13196 23024 13254
rect 17176 13010 19544 13080
rect 21052 13018 23024 13076
rect 17172 12838 19546 12896
rect 21052 12840 23024 12898
rect 17176 12654 19544 12724
rect 21052 12662 23024 12720
rect 17172 12482 19546 12540
rect 21052 12484 23024 12542
rect 17178 12298 19546 12368
rect 21052 12306 23024 12364
rect 17172 12126 19546 12184
rect 21052 12128 23024 12186
rect 17178 11942 19546 12012
rect 21052 11950 23024 12008
rect 17172 11770 19546 11828
rect 21052 11772 23024 11830
rect 17176 11586 19544 11656
rect 21052 11594 23024 11652
rect 17172 11414 19546 11472
rect 21052 11416 23024 11474
rect 17176 11230 19544 11300
rect 21052 11238 23024 11296
rect 17172 11058 19546 11116
rect 21052 11060 23024 11118
rect 17176 10874 19544 10944
rect 21052 10882 23024 10940
rect 17172 10702 19546 10760
rect 21052 10704 23024 10762
rect 17176 10518 19544 10588
rect 21052 10526 23024 10584
rect 17172 10346 19546 10404
rect 21052 10348 23024 10406
rect 17176 10162 19544 10232
rect 21052 10170 23024 10228
rect 17172 9990 19546 10048
rect 21052 9992 23024 10050
rect 17176 9806 19544 9876
rect 21052 9814 23024 9872
rect 17172 9634 19546 9692
rect 21052 9636 23024 9694
rect 17176 9450 19544 9520
rect 21052 9458 23024 9516
rect 17172 9278 19546 9336
rect 21052 9280 23024 9338
rect 17176 9094 19544 9164
rect 21052 9102 23024 9160
rect 17172 8922 19546 8980
rect 21052 8924 23024 8982
rect 17176 8738 19544 8808
rect 21052 8746 23024 8804
rect 17172 8566 19546 8624
rect 21052 8568 23024 8626
rect 17176 8382 19544 8452
rect 21054 8390 23026 8448
rect 17172 8210 19546 8268
rect 21052 8212 23024 8270
rect 17176 8026 19544 8096
rect 21052 8034 23024 8092
rect 17172 7854 19546 7912
rect 21052 7856 23024 7914
rect 17176 7670 19544 7740
rect 21052 7678 23024 7736
rect 17172 7498 19546 7556
rect 21052 7500 23024 7558
rect 17176 7314 19544 7384
rect 21052 7322 23024 7380
rect 17172 7140 19546 7198
rect 21052 7144 23024 7202
rect 17176 6958 19544 7028
rect 21052 6966 23024 7024
rect 17172 6786 19546 6844
rect 21052 6790 23024 6848
rect 17176 6602 19544 6672
rect 21052 6610 23024 6668
rect 17172 6430 19546 6488
rect 21052 6432 23024 6490
rect 17176 6246 19544 6316
rect 21052 6254 23024 6312
rect 17172 6074 19546 6132
rect 21052 6076 23024 6134
rect 17176 5890 19544 5960
rect 21052 5898 23024 5956
rect 17172 5718 19546 5776
rect 21052 5720 23024 5778
rect 17176 5534 19544 5604
rect 21052 5542 23024 5600
rect 17172 5362 19546 5420
rect 21052 5364 23024 5422
rect 17176 5178 19544 5248
rect 21052 5186 23024 5244
rect 17172 5006 19546 5064
rect 21052 5010 23024 5068
rect 17176 4822 19544 4892
rect 21052 4830 23024 4888
rect 17172 4650 19546 4708
rect 21052 4652 23024 4710
rect 17176 4466 19544 4536
rect 21052 4474 23024 4532
rect 17172 4294 19546 4352
rect 21052 4296 23024 4354
rect 17176 4110 19544 4180
rect 21052 4118 23024 4176
rect 17172 3936 19546 3994
rect 21052 3942 23024 4000
rect 17176 3754 19544 3824
rect 21052 3762 23024 3820
rect 17172 3582 19546 3640
rect 21052 3584 23024 3642
rect 17176 3398 19544 3468
rect 21052 3406 23024 3464
rect 17170 3226 19544 3284
rect 21052 3228 23024 3286
rect 17176 3042 19544 3112
rect 21052 3050 23024 3108
rect 17170 2870 19544 2928
rect 21052 2872 23024 2930
rect 25116 2734 25640 40588
rect 6242 1280 7252 2272
rect 11182 1294 12192 2286
rect 16524 1294 17534 2286
<< metal2 >>
rect 1996 38266 4954 44450
rect 23260 43860 27492 44454
rect 23260 43240 23738 43860
rect 27086 43240 27492 43860
rect 23260 41038 27492 43240
rect 23242 40588 27492 41038
rect 20646 40396 20656 40460
rect 23026 40396 23036 40460
rect 23242 40338 25116 40588
rect 20648 40280 20658 40338
rect 23028 40280 25116 40338
rect 20646 40160 20656 40224
rect 23026 40160 23036 40224
rect 20646 40046 20656 40104
rect 23026 40102 23036 40104
rect 23242 40102 25116 40280
rect 23026 40046 25116 40102
rect 20894 40044 25116 40046
rect 20644 39924 20654 39988
rect 23024 39924 23034 39988
rect 23242 39864 25116 40044
rect 20648 39806 20658 39864
rect 23028 39806 25116 39864
rect 20644 39688 20654 39752
rect 23024 39688 23034 39752
rect 23242 39632 25116 39806
rect 20646 39574 20656 39632
rect 23026 39574 25116 39632
rect 20646 39452 20656 39516
rect 23026 39452 23036 39516
rect 23242 39396 25116 39574
rect 20916 39394 25116 39396
rect 20646 39336 20656 39394
rect 23026 39338 25116 39394
rect 23026 39336 23036 39338
rect 20644 39214 20654 39278
rect 23024 39214 23034 39278
rect 20646 39102 20656 39160
rect 23026 39158 23036 39160
rect 23242 39158 25116 39338
rect 23026 39102 25116 39158
rect 20970 39100 25116 39102
rect 20646 38978 20656 39042
rect 23026 38978 23036 39042
rect 23242 38924 25116 39100
rect 20646 38866 20656 38924
rect 23026 38866 25116 38924
rect 20644 38746 20654 38810
rect 23024 38746 23034 38810
rect 23242 38688 25116 38866
rect 20894 38686 25116 38688
rect 20648 38628 20658 38686
rect 23028 38630 25116 38686
rect 23028 38628 23038 38630
rect 20646 38506 20656 38570
rect 23026 38506 23036 38570
rect 23242 38452 25116 38630
rect 20884 38450 25116 38452
rect 20646 38392 20656 38450
rect 23026 38394 25116 38450
rect 23026 38392 23036 38394
rect 20644 38270 20654 38334
rect 23024 38270 23034 38334
rect 1996 38084 2600 38266
rect 23242 38214 25116 38394
rect 3008 38138 3018 38204
rect 4792 38138 4802 38204
rect 20646 38156 20656 38214
rect 23026 38156 25116 38214
rect 1996 38080 3022 38084
rect 1996 38026 3012 38080
rect 4800 38026 4810 38080
rect 20644 38034 20654 38098
rect 23024 38034 23034 38098
rect 1996 37846 2600 38026
rect 23242 37980 25116 38156
rect 20922 37978 25116 37980
rect 3008 37902 3018 37968
rect 4792 37902 4802 37968
rect 20646 37920 20656 37978
rect 23026 37922 25116 37978
rect 23026 37920 23036 37922
rect 1996 37844 3026 37846
rect 1996 37790 3012 37844
rect 4800 37790 4810 37844
rect 20646 37798 20656 37862
rect 23026 37798 23036 37862
rect 1996 37788 3026 37790
rect 1996 37610 2600 37788
rect 23242 37744 25116 37922
rect 3008 37666 3018 37732
rect 4792 37666 4802 37732
rect 20648 37686 20658 37744
rect 23028 37686 25116 37744
rect 1996 37608 3024 37610
rect 1996 37554 3012 37608
rect 4800 37554 4810 37608
rect 20646 37562 20656 37626
rect 23026 37562 23036 37626
rect 1996 37552 3024 37554
rect 1996 37374 2600 37552
rect 23242 37506 25116 37686
rect 3008 37430 3018 37496
rect 4792 37430 4802 37496
rect 20646 37448 20656 37506
rect 23026 37448 25116 37506
rect 1996 37372 3030 37374
rect 1996 37318 3012 37372
rect 4800 37318 4810 37372
rect 20646 37326 20656 37390
rect 23026 37326 23036 37390
rect 1996 37316 3030 37318
rect 1996 37138 2600 37316
rect 23242 37272 25116 37448
rect 20906 37268 25116 37272
rect 3008 37194 3018 37260
rect 4792 37194 4802 37260
rect 20648 37210 20658 37268
rect 23028 37214 25116 37268
rect 23028 37210 23038 37214
rect 1996 37136 3022 37138
rect 1996 37082 3012 37136
rect 4800 37082 4810 37136
rect 20644 37092 20654 37156
rect 23024 37092 23034 37156
rect 1996 37080 3022 37082
rect 1996 36902 2600 37080
rect 23242 37036 25116 37214
rect 20932 37034 25116 37036
rect 3008 36958 3018 37024
rect 4792 36958 4802 37024
rect 20648 36976 20658 37034
rect 23028 36978 25116 37034
rect 23028 36976 23038 36978
rect 1996 36900 3028 36902
rect 1996 36846 3012 36900
rect 4800 36846 4810 36900
rect 20648 36856 20658 36920
rect 23028 36856 23038 36920
rect 1996 36844 3028 36846
rect 1996 36666 2600 36844
rect 23242 36798 25116 36978
rect 3008 36722 3018 36788
rect 4792 36722 4802 36788
rect 20648 36740 20658 36798
rect 23028 36740 25116 36798
rect 1996 36664 3022 36666
rect 1996 36610 3012 36664
rect 4800 36610 4810 36664
rect 20646 36618 20656 36682
rect 23026 36618 23036 36682
rect 1996 36608 3022 36610
rect 1996 36430 2600 36608
rect 3008 36486 3018 36552
rect 4792 36486 4802 36552
rect 20646 36504 20656 36562
rect 23026 36560 23036 36562
rect 23242 36560 25116 36740
rect 23026 36504 25116 36560
rect 20892 36502 25116 36504
rect 1996 36428 3026 36430
rect 1996 36374 3012 36428
rect 4800 36374 4810 36428
rect 20648 36382 20658 36446
rect 23028 36382 23038 36446
rect 1996 36372 3026 36374
rect 1996 36194 2600 36372
rect 23242 36328 25116 36502
rect 20884 36326 25116 36328
rect 3008 36250 3018 36316
rect 4792 36250 4802 36316
rect 20648 36268 20658 36326
rect 23028 36270 25116 36326
rect 23028 36268 23038 36270
rect 1996 36192 3028 36194
rect 1996 36138 3012 36192
rect 4800 36138 4810 36192
rect 20648 36146 20658 36210
rect 23028 36146 23038 36210
rect 1996 36136 3028 36138
rect 1996 35958 2600 36136
rect 23242 36092 25116 36270
rect 20920 36090 25116 36092
rect 3008 36014 3018 36080
rect 4792 36014 4802 36080
rect 20646 36032 20656 36090
rect 23026 36034 25116 36090
rect 23026 36032 23036 36034
rect 1996 35956 3044 35958
rect 1996 35902 3012 35956
rect 4800 35902 4810 35956
rect 20648 35912 20658 35976
rect 23028 35912 23038 35976
rect 1996 35900 3044 35902
rect 1996 35722 2600 35900
rect 3008 35778 3018 35844
rect 4792 35778 4802 35844
rect 20646 35798 20656 35856
rect 23026 35854 23036 35856
rect 23242 35854 25116 36034
rect 23026 35798 25116 35854
rect 20912 35796 25116 35798
rect 1996 35720 3034 35722
rect 1996 35666 3012 35720
rect 4800 35666 4810 35720
rect 20644 35674 20654 35738
rect 23024 35674 23034 35738
rect 1996 35664 3034 35666
rect 1996 35486 2600 35664
rect 23242 35620 25116 35796
rect 3008 35542 3018 35608
rect 4792 35542 4802 35608
rect 20648 35562 20658 35620
rect 23028 35562 25116 35620
rect 1996 35484 3048 35486
rect 1996 35430 3012 35484
rect 4800 35430 4810 35484
rect 20644 35436 20654 35500
rect 23024 35436 23034 35500
rect 1996 35428 3048 35430
rect 1996 35250 2600 35428
rect 23242 35384 25116 35562
rect 3008 35306 3018 35372
rect 4792 35306 4802 35372
rect 20646 35326 20656 35384
rect 23026 35326 25116 35384
rect 1996 35248 3038 35250
rect 1996 35194 3012 35248
rect 4800 35194 4810 35248
rect 20646 35202 20656 35266
rect 23026 35202 23036 35266
rect 1996 35192 3038 35194
rect 1996 35014 2600 35192
rect 23242 35148 25116 35326
rect 3008 35070 3018 35136
rect 4792 35070 4802 35136
rect 20646 35090 20656 35148
rect 23026 35090 25116 35148
rect 1996 35012 3052 35014
rect 1996 34958 3012 35012
rect 4800 34958 4810 35012
rect 20646 34966 20656 35030
rect 23026 34966 23036 35030
rect 1996 34956 3052 34958
rect 1996 34778 2600 34956
rect 23242 34910 25116 35090
rect 3008 34834 3018 34900
rect 4792 34834 4802 34900
rect 20646 34852 20656 34910
rect 23026 34852 25116 34910
rect 1996 34776 3052 34778
rect 1996 34722 3012 34776
rect 4800 34722 4810 34776
rect 20648 34730 20658 34794
rect 23028 34730 23038 34794
rect 1996 34720 3052 34722
rect 1996 34542 2600 34720
rect 23242 34676 25116 34852
rect 21004 34674 25116 34676
rect 3008 34598 3018 34664
rect 4792 34598 4802 34664
rect 20648 34616 20658 34674
rect 23028 34618 25116 34674
rect 23028 34616 23038 34618
rect 1996 34540 3056 34542
rect 1996 34486 3012 34540
rect 4800 34486 4810 34540
rect 20644 34496 20654 34560
rect 23024 34496 23034 34560
rect 1996 34484 3056 34486
rect 1996 34306 2600 34484
rect 23242 34440 25116 34618
rect 20942 34438 25116 34440
rect 3008 34362 3018 34428
rect 4792 34362 4802 34428
rect 20650 34380 20660 34438
rect 23030 34382 25116 34438
rect 23030 34380 23040 34382
rect 1996 34304 3048 34306
rect 1996 34250 3012 34304
rect 4800 34250 4810 34304
rect 20644 34258 20654 34322
rect 23024 34258 23034 34322
rect 1996 34248 3048 34250
rect 1996 34070 2600 34248
rect 23242 34202 25116 34382
rect 3008 34126 3018 34192
rect 4792 34126 4802 34192
rect 20648 34144 20658 34202
rect 23028 34144 25116 34202
rect 1996 34068 3032 34070
rect 1996 34014 3012 34068
rect 4800 34014 4810 34068
rect 20646 34024 20656 34088
rect 23026 34024 23036 34088
rect 1996 34012 3032 34014
rect 1996 33834 2600 34012
rect 23242 33966 25116 34144
rect 20900 33964 25116 33966
rect 3008 33890 3018 33956
rect 4792 33890 4802 33956
rect 20646 33906 20656 33964
rect 23026 33908 25116 33964
rect 23026 33906 23036 33908
rect 1996 33832 3026 33834
rect 1996 33778 3012 33832
rect 4800 33778 4810 33832
rect 20646 33786 20656 33850
rect 23026 33786 23036 33850
rect 1996 33776 3026 33778
rect 1996 33598 2600 33776
rect 23242 33732 25116 33908
rect 3008 33654 3018 33720
rect 4792 33654 4802 33720
rect 20646 33674 20656 33732
rect 23026 33674 25116 33732
rect 1996 33596 3042 33598
rect 1996 33542 3012 33596
rect 4800 33542 4810 33596
rect 20646 33550 20656 33614
rect 23026 33550 23036 33614
rect 1996 33540 3042 33542
rect 1996 33362 2600 33540
rect 23242 33494 25116 33674
rect 3008 33418 3018 33484
rect 4792 33418 4802 33484
rect 20646 33436 20656 33494
rect 23026 33436 25116 33494
rect 1996 33360 3046 33362
rect 1996 33306 3012 33360
rect 4800 33306 4810 33360
rect 20646 33316 20656 33380
rect 23026 33316 23036 33380
rect 1996 33304 3046 33306
rect 1996 33126 2600 33304
rect 3008 33182 3018 33248
rect 4792 33182 4802 33248
rect 20648 33202 20658 33260
rect 23028 33258 23038 33260
rect 23242 33258 25116 33436
rect 23028 33202 25116 33258
rect 20900 33200 25116 33202
rect 1996 33124 3054 33126
rect 1996 33070 3012 33124
rect 4800 33070 4810 33124
rect 20646 33080 20656 33144
rect 23026 33080 23036 33144
rect 1996 33068 3054 33070
rect 1996 32890 2600 33068
rect 23242 33024 25116 33200
rect 20894 33022 25116 33024
rect 3008 32946 3018 33012
rect 4792 32946 4802 33012
rect 20648 32964 20658 33022
rect 23028 32966 25116 33022
rect 23028 32964 23038 32966
rect 1996 32888 3058 32890
rect 1996 32834 3012 32888
rect 4800 32834 4810 32888
rect 20646 32842 20656 32906
rect 23026 32842 23036 32906
rect 1996 32832 3058 32834
rect 1996 32656 2600 32832
rect 23242 32788 25116 32966
rect 3008 32710 3018 32776
rect 4792 32710 4802 32776
rect 20646 32730 20656 32788
rect 23026 32730 25116 32788
rect 1996 32652 3034 32656
rect 1996 32598 3012 32652
rect 4800 32598 4810 32652
rect 20648 32608 20658 32672
rect 23028 32608 23038 32672
rect 1996 32418 2600 32598
rect 3008 32474 3018 32540
rect 4792 32474 4802 32540
rect 20646 32494 20656 32552
rect 23026 32550 23036 32552
rect 23242 32550 25116 32730
rect 23026 32494 25116 32550
rect 20936 32492 25116 32494
rect 1996 32416 3034 32418
rect 1996 32362 3012 32416
rect 4800 32362 4810 32416
rect 20648 32374 20658 32438
rect 23028 32374 23038 32438
rect 1996 32360 3034 32362
rect 1996 32182 2600 32360
rect 23242 32314 25116 32492
rect 3008 32238 3018 32304
rect 4792 32238 4802 32304
rect 20646 32256 20656 32314
rect 23026 32256 25116 32314
rect 1996 32180 3022 32182
rect 1996 32126 3012 32180
rect 4800 32126 4810 32180
rect 20646 32134 20656 32198
rect 23026 32134 23036 32198
rect 1996 32124 3022 32126
rect 1996 31946 2600 32124
rect 23242 32078 25116 32256
rect 3008 32002 3018 32068
rect 4792 32002 4802 32068
rect 20646 32020 20656 32078
rect 23026 32020 25116 32078
rect 1996 31944 3056 31946
rect 1996 31890 3012 31944
rect 4800 31890 4810 31944
rect 20646 31900 20656 31964
rect 23026 31900 23036 31964
rect 1996 31888 3056 31890
rect 1996 31710 2600 31888
rect 23242 31840 25116 32020
rect 3006 31766 3016 31832
rect 4790 31766 4800 31832
rect 20648 31782 20658 31840
rect 23028 31782 25116 31840
rect 1996 31708 3022 31710
rect 1996 31654 3012 31708
rect 4800 31654 4810 31708
rect 20646 31662 20656 31726
rect 23026 31662 23036 31726
rect 1996 31652 3022 31654
rect 1996 31474 2600 31652
rect 23242 31606 25116 31782
rect 3008 31530 3018 31596
rect 4792 31530 4802 31596
rect 20648 31548 20658 31606
rect 23028 31548 25116 31606
rect 1996 31472 3066 31474
rect 1996 31418 3012 31472
rect 4800 31418 4810 31472
rect 20646 31428 20656 31492
rect 23026 31428 23036 31492
rect 1996 31416 3066 31418
rect 1996 31238 2600 31416
rect 23242 31372 25116 31548
rect 3008 31294 3018 31360
rect 4792 31294 4802 31360
rect 20648 31314 20658 31372
rect 23028 31314 25116 31372
rect 1996 31236 3032 31238
rect 1996 31182 3012 31236
rect 4800 31182 4810 31236
rect 20646 31192 20656 31256
rect 23026 31192 23036 31256
rect 1996 31180 3032 31182
rect 1996 30994 2600 31180
rect 23242 31136 25116 31314
rect 20900 31134 25116 31136
rect 3008 31060 3018 31120
rect 4792 31060 4802 31120
rect 20646 31076 20656 31134
rect 23026 31078 25116 31134
rect 23026 31076 23036 31078
rect 1996 30836 4398 30994
rect 20644 30956 20654 31020
rect 23024 30956 23034 31020
rect 20646 30842 20656 30900
rect 23026 30898 23036 30900
rect 23242 30898 25116 31078
rect 23026 30842 25116 30898
rect 20884 30840 25116 30842
rect 1996 29890 4400 30836
rect 20646 30718 20656 30782
rect 23026 30718 23036 30782
rect 23242 30662 25116 30840
rect 20646 30604 20656 30662
rect 23026 30604 25116 30662
rect 20646 30482 20656 30546
rect 23026 30482 23036 30546
rect 23242 30426 25116 30604
rect 20646 30368 20656 30426
rect 23026 30368 25116 30426
rect 20646 30248 20656 30312
rect 23026 30248 23036 30312
rect 23242 30190 25116 30368
rect 21062 30188 25116 30190
rect 20648 30130 20658 30188
rect 23028 30132 25116 30188
rect 23028 30130 23038 30132
rect 20646 30010 20656 30074
rect 23026 30010 23036 30074
rect 23242 29954 25116 30132
rect 20648 29896 20658 29954
rect 23028 29896 25116 29954
rect 1996 3110 2784 29890
rect 3772 15586 4400 29890
rect 20648 29776 20658 29840
rect 23028 29776 23038 29840
rect 23242 27192 25116 29896
rect 20430 25230 20756 25298
rect 20904 25230 21006 25240
rect 20430 25226 23024 25230
rect 20430 25170 21052 25226
rect 23024 25170 23034 25226
rect 20430 25168 23024 25170
rect 20430 24876 20756 25168
rect 20904 24876 20926 25168
rect 20430 24814 20926 24876
rect 20430 24520 20756 24814
rect 20904 24520 20926 24814
rect 20430 24458 20926 24520
rect 20430 24164 20756 24458
rect 20904 24164 20926 24458
rect 20430 24102 20926 24164
rect 20430 23808 20756 24102
rect 20904 23808 20926 24102
rect 20430 23746 20926 23808
rect 20430 23452 20756 23746
rect 20904 23452 20926 23746
rect 20430 23390 20926 23452
rect 20430 23096 20756 23390
rect 20904 23096 20926 23390
rect 20430 23034 20926 23096
rect 20430 23032 20756 23034
rect 19814 22772 19974 22782
rect 18478 22684 18982 22694
rect 19814 22650 19974 22660
rect 20432 22740 20756 23032
rect 20904 22740 20926 23034
rect 20432 22678 20926 22740
rect 18478 22284 18982 22294
rect 20432 22384 20756 22678
rect 20904 22384 20926 22678
rect 20432 22322 20926 22384
rect 7996 22038 8448 22044
rect 20432 22038 20756 22322
rect 7996 21218 20756 22038
rect 7996 20730 8448 21218
rect 19810 21144 19970 21154
rect 19788 21030 19810 21144
rect 19970 21030 20220 21144
rect 19810 21020 19970 21030
rect 20010 20832 20220 21030
rect 20430 20960 20756 21218
rect 20904 20960 20926 22322
rect 20430 20898 20926 20960
rect 7996 20666 9172 20730
rect 11542 20666 11808 20730
rect 14178 20666 14188 20730
rect 19950 20728 20276 20832
rect 14526 20670 14536 20728
rect 16910 20670 17172 20728
rect 19546 20670 20276 20728
rect 7996 20374 8448 20666
rect 9162 20486 9172 20556
rect 11542 20486 11552 20556
rect 11798 20486 11808 20556
rect 14176 20486 14186 20556
rect 14530 20488 14540 20558
rect 16908 20488 16918 20558
rect 17166 20486 17176 20556
rect 19544 20486 19554 20556
rect 7996 20310 9172 20374
rect 11542 20310 11808 20374
rect 14178 20310 14188 20374
rect 19950 20372 20276 20670
rect 14526 20314 14536 20372
rect 16910 20314 17172 20372
rect 19546 20314 20276 20372
rect 7996 20018 8448 20310
rect 9162 20130 9172 20200
rect 11540 20130 11550 20200
rect 11798 20130 11808 20200
rect 14176 20130 14186 20200
rect 14530 20130 14540 20200
rect 16908 20130 16918 20200
rect 17166 20130 17176 20200
rect 19544 20130 19554 20200
rect 19950 20018 20276 20314
rect 7996 19954 9172 20018
rect 11542 19954 11808 20018
rect 14178 19954 14188 20018
rect 17606 20016 20276 20018
rect 14526 19958 14536 20016
rect 16910 19958 17172 20016
rect 19546 19960 20276 20016
rect 19546 19958 19556 19960
rect 7996 19662 8448 19954
rect 9162 19774 9172 19844
rect 11540 19774 11550 19844
rect 11798 19774 11808 19844
rect 14176 19774 14186 19844
rect 14530 19774 14540 19844
rect 16908 19774 16918 19844
rect 17166 19774 17176 19844
rect 19544 19774 19554 19844
rect 7996 19598 9172 19662
rect 11542 19598 11808 19662
rect 14178 19598 14188 19662
rect 14526 19602 14536 19660
rect 16910 19602 17172 19660
rect 19546 19658 19556 19660
rect 19950 19658 20276 19960
rect 19546 19602 20276 19658
rect 17598 19600 20276 19602
rect 7996 19308 8448 19598
rect 9162 19420 9172 19490
rect 11540 19420 11550 19490
rect 11798 19418 11808 19488
rect 14176 19418 14186 19488
rect 14530 19416 14540 19486
rect 16908 19416 16918 19486
rect 17166 19416 17176 19486
rect 19544 19416 19554 19486
rect 7996 19244 9172 19308
rect 11542 19244 11808 19308
rect 14178 19244 14188 19308
rect 19950 19304 20276 19600
rect 14526 19246 14536 19304
rect 16910 19246 17172 19304
rect 19546 19246 20276 19304
rect 7996 18950 8448 19244
rect 9162 19062 9172 19132
rect 11540 19062 11550 19132
rect 11798 19062 11808 19132
rect 14176 19062 14186 19132
rect 14530 19062 14540 19132
rect 16908 19062 16918 19132
rect 17166 19062 17176 19132
rect 19544 19062 19554 19132
rect 7996 18886 9172 18950
rect 11542 18886 11808 18950
rect 14178 18886 14188 18950
rect 19950 18948 20276 19246
rect 14526 18890 14536 18948
rect 16910 18890 17172 18948
rect 19546 18890 20276 18948
rect 7996 18594 8448 18886
rect 9162 18706 9172 18776
rect 11540 18706 11550 18776
rect 11798 18706 11808 18776
rect 14176 18706 14186 18776
rect 14530 18706 14540 18776
rect 16908 18706 16918 18776
rect 17166 18706 17176 18776
rect 19544 18706 19554 18776
rect 7996 18530 9172 18594
rect 11542 18530 11808 18594
rect 14178 18530 14188 18594
rect 19950 18592 20276 18890
rect 14526 18534 14536 18592
rect 16910 18534 17172 18592
rect 19546 18534 20276 18592
rect 7996 18238 8448 18530
rect 9162 18350 9172 18420
rect 11540 18350 11550 18420
rect 11798 18350 11808 18420
rect 14176 18350 14186 18420
rect 14530 18350 14540 18420
rect 16908 18350 16918 18420
rect 17166 18350 17176 18420
rect 19544 18350 19554 18420
rect 19950 18238 20276 18534
rect 7996 18174 9172 18238
rect 11542 18174 11808 18238
rect 14178 18174 14188 18238
rect 17608 18236 20276 18238
rect 14526 18178 14536 18236
rect 16910 18178 17172 18236
rect 19546 18180 20276 18236
rect 19546 18178 19556 18180
rect 7996 17882 8448 18174
rect 9162 17994 9172 18064
rect 11540 17994 11550 18064
rect 11798 17994 11808 18064
rect 14176 17994 14186 18064
rect 14530 17994 14540 18064
rect 16908 17994 16918 18064
rect 17166 17994 17176 18064
rect 19544 17994 19554 18064
rect 7996 17818 9172 17882
rect 11542 17818 11808 17882
rect 14178 17818 14188 17882
rect 19950 17880 20276 18180
rect 14526 17822 14536 17880
rect 16910 17822 17172 17880
rect 19546 17822 20276 17880
rect 7996 17528 8448 17818
rect 9162 17638 9172 17708
rect 11540 17638 11550 17708
rect 11798 17638 11808 17708
rect 14176 17638 14186 17708
rect 14530 17638 14540 17708
rect 16908 17638 16918 17708
rect 17166 17636 17176 17706
rect 19544 17636 19554 17706
rect 7996 17464 9172 17528
rect 11542 17464 11808 17528
rect 14178 17464 14188 17528
rect 19950 17524 20276 17822
rect 14526 17466 14536 17524
rect 16910 17466 17172 17524
rect 19546 17466 20276 17524
rect 7996 17172 8448 17464
rect 9162 17280 9172 17352
rect 11540 17280 11550 17352
rect 11798 17282 11808 17352
rect 14176 17282 14186 17352
rect 14530 17282 14540 17352
rect 16908 17282 16918 17352
rect 17166 17282 17176 17352
rect 19544 17282 19554 17352
rect 7996 17108 9172 17172
rect 11542 17108 11808 17172
rect 14178 17108 14188 17172
rect 19950 17168 20276 17466
rect 14526 17110 14536 17168
rect 16910 17110 17172 17168
rect 19546 17110 20276 17168
rect 7996 16816 8448 17108
rect 9162 16926 9172 16996
rect 11540 16926 11550 16996
rect 11798 16926 11808 16996
rect 14176 16926 14186 16996
rect 14530 16926 14540 16996
rect 16908 16926 16918 16996
rect 17166 16926 17176 16996
rect 19544 16926 19554 16996
rect 7996 16752 9172 16816
rect 11542 16752 11808 16816
rect 14178 16752 14188 16816
rect 19950 16812 20276 17110
rect 14526 16754 14536 16812
rect 16910 16754 17172 16812
rect 19546 16754 20276 16812
rect 7996 16460 8448 16752
rect 9162 16570 9172 16640
rect 11540 16570 11550 16640
rect 11798 16570 11808 16640
rect 14176 16570 14186 16640
rect 14530 16570 14540 16640
rect 16908 16570 16918 16640
rect 17166 16570 17176 16640
rect 19544 16570 19554 16640
rect 9162 16460 9172 16462
rect 7996 16398 9172 16460
rect 11542 16460 11552 16462
rect 11542 16398 11808 16460
rect 7996 16396 11808 16398
rect 14178 16396 14188 16460
rect 19950 16458 20276 16754
rect 17606 16456 20276 16458
rect 14526 16398 14536 16456
rect 16910 16398 17172 16456
rect 19546 16400 20276 16456
rect 19546 16398 19556 16400
rect 7996 16102 8448 16396
rect 9162 16214 9172 16286
rect 11540 16214 11550 16286
rect 11798 16216 11808 16286
rect 14176 16216 14186 16286
rect 14530 16214 14540 16284
rect 16908 16214 16918 16284
rect 17166 16214 17176 16284
rect 19544 16214 19554 16284
rect 7996 16038 9172 16102
rect 11542 16038 11808 16102
rect 14178 16038 14188 16102
rect 19950 16100 20276 16400
rect 14526 16042 14536 16100
rect 16910 16042 17172 16100
rect 19546 16042 20276 16100
rect 7996 15746 8448 16038
rect 9162 15858 9172 15928
rect 11540 15858 11550 15928
rect 11798 15858 11808 15928
rect 14176 15858 14186 15928
rect 14530 15856 14540 15926
rect 16908 15856 16918 15926
rect 17166 15858 17176 15928
rect 19544 15858 19554 15928
rect 19950 15746 20276 16042
rect 4770 15648 4780 15710
rect 6568 15648 6578 15710
rect 7996 15682 9172 15746
rect 11542 15682 11808 15746
rect 14178 15682 14188 15746
rect 17628 15744 20276 15746
rect 14526 15686 14536 15744
rect 16910 15686 17172 15744
rect 19546 15688 20276 15744
rect 19546 15686 19556 15688
rect 4772 15586 4782 15588
rect 3772 15536 4782 15586
rect 3772 15350 4398 15536
rect 4772 15534 4782 15536
rect 6570 15534 6580 15588
rect 4770 15412 4780 15474
rect 6568 15412 6578 15474
rect 7996 15392 8448 15682
rect 9162 15502 9172 15572
rect 11540 15502 11550 15572
rect 11798 15502 11808 15572
rect 14176 15502 14186 15572
rect 14530 15502 14540 15572
rect 16908 15502 16918 15572
rect 17166 15502 17176 15572
rect 19544 15502 19554 15572
rect 4772 15350 4782 15352
rect 3772 15300 4782 15350
rect 3772 15114 4398 15300
rect 4772 15298 4782 15300
rect 6570 15298 6580 15352
rect 7996 15328 9172 15392
rect 11542 15328 11808 15392
rect 14178 15328 14188 15392
rect 19950 15388 20276 15688
rect 14526 15330 14536 15388
rect 16910 15330 17172 15388
rect 19546 15330 20276 15388
rect 4770 15176 4780 15238
rect 6568 15176 6578 15238
rect 4772 15114 4782 15116
rect 3772 15064 4782 15114
rect 3772 14878 4398 15064
rect 4772 15062 4782 15064
rect 6570 15062 6580 15116
rect 7996 15034 8448 15328
rect 9162 15146 9172 15216
rect 11540 15146 11550 15216
rect 11798 15146 11808 15216
rect 14176 15146 14186 15216
rect 14530 15146 14540 15216
rect 16908 15146 16918 15216
rect 17166 15146 17176 15216
rect 19544 15146 19554 15216
rect 4770 14940 4780 15002
rect 6568 14940 6578 15002
rect 7996 14970 9172 15034
rect 11542 14970 11808 15034
rect 14178 14970 14188 15034
rect 19950 15032 20276 15330
rect 14526 14974 14536 15032
rect 16910 14974 17172 15032
rect 19546 14974 20276 15032
rect 4772 14878 4782 14880
rect 3772 14828 4782 14878
rect 3772 14642 4398 14828
rect 4772 14826 4782 14828
rect 6570 14826 6580 14880
rect 4770 14704 4780 14766
rect 6568 14704 6578 14766
rect 7996 14680 8448 14970
rect 9162 14790 9172 14860
rect 11540 14790 11550 14860
rect 11798 14790 11808 14860
rect 14176 14790 14186 14860
rect 14530 14790 14540 14860
rect 16908 14790 16918 14860
rect 17166 14790 17176 14860
rect 19544 14790 19554 14860
rect 4772 14642 4782 14644
rect 3772 14592 4782 14642
rect 3772 14408 4398 14592
rect 4772 14590 4782 14592
rect 6570 14590 6580 14644
rect 7996 14616 9172 14680
rect 11542 14616 11808 14680
rect 14178 14616 14188 14680
rect 19950 14678 20276 14974
rect 17596 14676 20276 14678
rect 14526 14618 14536 14676
rect 16910 14618 17172 14676
rect 19546 14620 20276 14676
rect 19546 14618 19556 14620
rect 4770 14468 4780 14530
rect 6568 14468 6578 14530
rect 3772 14358 4782 14408
rect 3772 14170 4398 14358
rect 4772 14354 4782 14358
rect 6570 14354 6580 14408
rect 7996 14322 8448 14616
rect 9162 14434 9172 14504
rect 11540 14434 11550 14504
rect 11798 14434 11808 14504
rect 14176 14434 14186 14504
rect 14530 14434 14540 14504
rect 16908 14434 16918 14504
rect 17166 14434 17176 14504
rect 19544 14434 19554 14504
rect 4770 14232 4780 14294
rect 6568 14232 6578 14294
rect 7996 14258 9172 14322
rect 11542 14258 11808 14322
rect 14178 14258 14188 14322
rect 14526 14262 14536 14320
rect 16910 14318 19546 14320
rect 19950 14318 20276 14620
rect 16910 14262 17172 14318
rect 17162 14260 17172 14262
rect 19546 14260 20276 14318
rect 4770 14170 4780 14172
rect 3772 14120 4780 14170
rect 3772 13934 4398 14120
rect 4770 14118 4780 14120
rect 6568 14118 6578 14172
rect 4768 13996 4778 14058
rect 6568 13996 6578 14058
rect 7996 13968 8448 14258
rect 9162 14078 9172 14148
rect 11540 14078 11550 14148
rect 11798 14078 11808 14148
rect 14176 14078 14186 14148
rect 14530 14076 14540 14146
rect 16908 14076 16918 14146
rect 17166 14078 17176 14148
rect 19544 14078 19554 14148
rect 19950 13968 20276 14260
rect 20430 20604 20756 20898
rect 20904 20604 20926 20898
rect 20430 20542 20926 20604
rect 20430 20248 20756 20542
rect 20904 20248 20926 20542
rect 20430 20186 20926 20248
rect 20430 19892 20756 20186
rect 20904 19892 20926 20186
rect 20430 19830 20926 19892
rect 20430 19536 20756 19830
rect 20904 19536 20926 19830
rect 20430 19474 20926 19536
rect 20430 19180 20756 19474
rect 20904 19180 20926 19474
rect 20430 19118 20926 19180
rect 20430 18824 20756 19118
rect 20904 18824 20926 19118
rect 20430 18762 20926 18824
rect 20430 18468 20756 18762
rect 20904 18468 20926 18762
rect 20430 18406 20926 18468
rect 20430 18112 20756 18406
rect 20904 18112 20926 18406
rect 20430 18050 20926 18112
rect 20430 17756 20756 18050
rect 20904 17756 20926 18050
rect 20430 17694 20926 17756
rect 20430 17400 20756 17694
rect 20904 17400 20926 17694
rect 20430 17338 20926 17400
rect 20430 17044 20756 17338
rect 20904 17044 20926 17338
rect 20430 16982 20926 17044
rect 20430 16688 20756 16982
rect 20904 16688 20926 16982
rect 20430 16626 20926 16688
rect 20430 16332 20756 16626
rect 20904 16332 20926 16626
rect 20430 16270 20926 16332
rect 20430 15976 20756 16270
rect 20904 15976 20926 16270
rect 20430 15914 20926 15976
rect 20430 15620 20756 15914
rect 20904 15620 20926 15914
rect 20430 15558 20926 15620
rect 20430 15264 20756 15558
rect 20904 15264 20926 15558
rect 20430 15202 20926 15264
rect 20430 14908 20756 15202
rect 20904 14908 20926 15202
rect 20430 14846 20926 14908
rect 20430 14552 20756 14846
rect 20904 14552 20926 14846
rect 20430 14490 20926 14552
rect 20430 14194 20756 14490
rect 20904 14194 20926 14490
rect 21000 24876 21006 25168
rect 21044 24992 21054 25056
rect 23024 24992 23034 25056
rect 21000 24872 23024 24876
rect 21000 24816 21052 24872
rect 23024 24816 23034 24872
rect 21000 24814 23024 24816
rect 21000 24520 21006 24814
rect 21044 24636 21054 24700
rect 23024 24636 23034 24700
rect 21000 24516 23024 24520
rect 21000 24460 21052 24516
rect 23024 24460 23034 24516
rect 21000 24458 23024 24460
rect 21000 24164 21006 24458
rect 21044 24278 21054 24342
rect 23024 24278 23034 24342
rect 21000 24160 23024 24164
rect 21000 24104 21052 24160
rect 23024 24104 23034 24160
rect 21000 24102 23024 24104
rect 21000 23808 21006 24102
rect 21044 23922 21054 23986
rect 23024 23922 23034 23986
rect 21000 23804 23024 23808
rect 21000 23748 21052 23804
rect 23024 23748 23034 23804
rect 21000 23746 23024 23748
rect 21000 23452 21006 23746
rect 21042 23568 21052 23632
rect 23022 23568 23032 23632
rect 21000 23448 23024 23452
rect 21000 23392 21052 23448
rect 23024 23392 23034 23448
rect 21000 23390 23024 23392
rect 21000 23096 21006 23390
rect 21044 23210 21054 23274
rect 23024 23210 23034 23274
rect 21000 23092 23024 23096
rect 21000 23036 21052 23092
rect 23024 23036 23034 23092
rect 21000 23034 23024 23036
rect 21000 22740 21006 23034
rect 21044 22856 21054 22920
rect 23024 22856 23034 22920
rect 21000 22736 23024 22740
rect 21000 22680 21052 22736
rect 23024 22680 23034 22736
rect 21000 22678 23024 22680
rect 21000 22384 21006 22678
rect 21044 22498 21054 22562
rect 23024 22498 23034 22562
rect 21000 22380 23024 22384
rect 21000 22324 21052 22380
rect 23024 22324 23034 22380
rect 21000 22322 23024 22324
rect 21000 22028 21006 22322
rect 21044 22142 21054 22206
rect 23024 22142 23034 22206
rect 21000 22024 23024 22028
rect 21000 21968 21052 22024
rect 23024 21968 23034 22024
rect 21000 21966 23024 21968
rect 21000 21672 21006 21966
rect 21044 21788 21054 21852
rect 23024 21788 23034 21852
rect 21000 21668 23024 21672
rect 21000 21612 21052 21668
rect 23024 21612 23034 21668
rect 21000 21610 23024 21612
rect 21000 21316 21006 21610
rect 21044 21430 21054 21494
rect 23024 21430 23034 21494
rect 21000 21312 23020 21316
rect 21000 21256 21052 21312
rect 23024 21256 23034 21312
rect 21000 21254 23020 21256
rect 21000 20960 21006 21254
rect 21044 21076 21054 21140
rect 23024 21076 23034 21140
rect 21000 20956 23024 20960
rect 21000 20900 21052 20956
rect 23024 20900 23034 20956
rect 21000 20898 23024 20900
rect 21000 20604 21006 20898
rect 21042 20718 21052 20782
rect 23022 20718 23032 20782
rect 21000 20600 23024 20604
rect 21000 20544 21052 20600
rect 23024 20544 23034 20600
rect 21000 20542 23024 20544
rect 21000 20248 21006 20542
rect 21044 20360 21054 20424
rect 23024 20360 23034 20424
rect 21000 20244 23024 20248
rect 21000 20188 21052 20244
rect 23024 20188 23034 20244
rect 21000 20186 23024 20188
rect 21000 19892 21006 20186
rect 21042 20008 21052 20072
rect 23022 20008 23032 20072
rect 21000 19888 23024 19892
rect 21000 19832 21052 19888
rect 23024 19832 23034 19888
rect 21000 19830 23024 19832
rect 21000 19536 21006 19830
rect 21044 19650 21054 19714
rect 23024 19650 23034 19714
rect 21000 19532 23024 19536
rect 21000 19476 21052 19532
rect 23024 19476 23034 19532
rect 21000 19474 23024 19476
rect 21000 19180 21006 19474
rect 21042 19296 21052 19360
rect 23022 19296 23032 19360
rect 21000 19176 23024 19180
rect 21000 19120 21052 19176
rect 23024 19120 23034 19176
rect 21000 19118 23024 19120
rect 21000 18824 21006 19118
rect 21044 18938 21054 19002
rect 23024 18938 23034 19002
rect 21000 18820 23024 18824
rect 21000 18764 21052 18820
rect 23024 18764 23034 18820
rect 21000 18762 23024 18764
rect 21000 18468 21006 18762
rect 21042 18582 21052 18646
rect 23022 18582 23032 18646
rect 21000 18464 23024 18468
rect 21000 18408 21052 18464
rect 23024 18408 23034 18464
rect 21000 18406 23024 18408
rect 21000 18112 21006 18406
rect 21044 18226 21054 18290
rect 23024 18226 23034 18290
rect 21000 18108 23024 18112
rect 21000 18052 21052 18108
rect 23024 18052 23034 18108
rect 21000 18050 23024 18052
rect 21000 17756 21006 18050
rect 21044 17870 21054 17934
rect 23024 17870 23034 17934
rect 21000 17752 23024 17756
rect 21000 17696 21052 17752
rect 23024 17696 23034 17752
rect 21000 17694 23024 17696
rect 21000 17400 21006 17694
rect 21044 17514 21054 17578
rect 23024 17514 23034 17578
rect 21000 17396 23024 17400
rect 21000 17340 21052 17396
rect 23024 17340 23034 17396
rect 21000 17338 23024 17340
rect 21000 17044 21006 17338
rect 21044 17158 21054 17222
rect 23024 17158 23034 17222
rect 21000 17040 23024 17044
rect 21000 16984 21052 17040
rect 23024 16984 23034 17040
rect 21000 16982 23024 16984
rect 21000 16688 21006 16982
rect 21044 16802 21054 16866
rect 23024 16802 23034 16866
rect 21000 16684 23024 16688
rect 21000 16628 21052 16684
rect 23024 16628 23034 16684
rect 21000 16626 23024 16628
rect 21000 16332 21006 16626
rect 21042 16446 21052 16510
rect 23022 16446 23032 16510
rect 21000 16328 23024 16332
rect 21000 16272 21052 16328
rect 23024 16272 23034 16328
rect 21000 16270 23024 16272
rect 21000 15976 21006 16270
rect 21044 16090 21054 16154
rect 23024 16090 23034 16154
rect 21000 15972 23024 15976
rect 21000 15916 21052 15972
rect 23024 15916 23034 15972
rect 21000 15914 23024 15916
rect 21000 15620 21006 15914
rect 21044 15736 21054 15800
rect 23024 15736 23034 15800
rect 21000 15616 23024 15620
rect 21000 15560 21052 15616
rect 23024 15560 23034 15616
rect 21000 15558 23024 15560
rect 21000 15264 21006 15558
rect 21044 15378 21054 15442
rect 23024 15378 23034 15442
rect 21000 15260 23024 15264
rect 21000 15204 21052 15260
rect 23024 15204 23034 15260
rect 21000 15202 23024 15204
rect 21000 14908 21006 15202
rect 21044 15022 21054 15086
rect 23024 15022 23034 15086
rect 21000 14904 23024 14908
rect 21000 14848 21052 14904
rect 23024 14848 23034 14904
rect 21000 14846 23024 14848
rect 21000 14552 21006 14846
rect 21044 14668 21054 14732
rect 23024 14668 23034 14732
rect 21000 14548 23024 14552
rect 21000 14492 21052 14548
rect 23024 14492 23034 14548
rect 21000 14490 23024 14492
rect 21000 14194 21006 14490
rect 21044 14310 21054 14374
rect 23024 14310 23034 14374
rect 20430 14192 23024 14194
rect 20430 14136 21052 14192
rect 23024 14136 23034 14192
rect 20430 14134 23024 14136
rect 20430 14098 20756 14134
rect 20904 14132 21006 14134
rect 4770 13934 4780 13936
rect 3772 13884 4780 13934
rect 3772 13698 4398 13884
rect 4770 13882 4780 13884
rect 6568 13882 6578 13936
rect 7996 13904 9172 13968
rect 11542 13904 11808 13968
rect 14178 13904 14188 13968
rect 14526 13906 14536 13964
rect 16910 13906 17172 13964
rect 19546 13962 19556 13964
rect 19950 13962 21052 13968
rect 19546 13910 21052 13962
rect 23024 13910 23034 13968
rect 19546 13908 23024 13910
rect 19546 13906 20276 13908
rect 17606 13904 20276 13906
rect 4770 13760 4780 13822
rect 6568 13760 6578 13822
rect 4772 13698 4782 13700
rect 3772 13648 4782 13698
rect 3772 13462 4398 13648
rect 4772 13646 4782 13648
rect 6570 13646 6580 13700
rect 7996 13612 8448 13904
rect 9162 13722 9172 13792
rect 11540 13722 11550 13792
rect 11798 13722 11808 13792
rect 14176 13722 14186 13792
rect 14530 13722 14540 13792
rect 16908 13722 16918 13792
rect 17166 13722 17176 13792
rect 19544 13722 19554 13792
rect 9162 13612 9172 13614
rect 4770 13524 4780 13586
rect 6568 13524 6578 13586
rect 7996 13550 9172 13612
rect 11542 13612 11552 13614
rect 11542 13550 11808 13612
rect 7996 13548 11808 13550
rect 14178 13548 14188 13612
rect 19950 13610 20276 13904
rect 20594 13610 21008 13908
rect 21042 13730 21052 13788
rect 23024 13730 23034 13788
rect 19950 13608 21052 13610
rect 14526 13550 14536 13608
rect 16910 13550 17172 13608
rect 19546 13552 21052 13608
rect 23024 13552 23034 13610
rect 19546 13550 23020 13552
rect 4772 13462 4782 13464
rect 3772 13412 4782 13462
rect 3772 13226 4398 13412
rect 4772 13410 4782 13412
rect 6570 13410 6580 13464
rect 4770 13288 4780 13350
rect 6568 13288 6578 13350
rect 7996 13254 8448 13548
rect 9162 13366 9172 13436
rect 11540 13366 11550 13436
rect 11798 13366 11808 13436
rect 14176 13366 14186 13436
rect 14530 13366 14540 13436
rect 16908 13366 16918 13436
rect 17166 13366 17176 13436
rect 19544 13366 19554 13436
rect 9162 13254 9172 13256
rect 4772 13226 4782 13228
rect 3772 13176 4782 13226
rect 3772 12990 4398 13176
rect 4772 13174 4782 13176
rect 6570 13174 6580 13228
rect 7996 13192 9172 13254
rect 11542 13254 11552 13256
rect 19950 13254 20276 13550
rect 20594 13254 21008 13550
rect 21042 13374 21052 13432
rect 23024 13374 23034 13432
rect 11542 13192 11808 13254
rect 7996 13190 11808 13192
rect 14178 13190 14188 13254
rect 14526 13194 14536 13252
rect 16910 13194 17172 13252
rect 19546 13250 19556 13252
rect 19950 13250 21052 13254
rect 19546 13196 21052 13250
rect 23024 13196 23034 13254
rect 19546 13194 23024 13196
rect 17648 13192 20276 13194
rect 4770 13052 4780 13114
rect 6568 13052 6578 13114
rect 4772 12990 4782 12992
rect 3772 12940 4782 12990
rect 3772 12754 4398 12940
rect 4772 12938 4782 12940
rect 6570 12938 6580 12992
rect 7996 12898 8448 13190
rect 9162 13010 9172 13080
rect 11540 13010 11550 13080
rect 11798 13010 11808 13080
rect 14176 13010 14186 13080
rect 14530 13010 14540 13080
rect 16908 13010 16918 13080
rect 17166 13010 17176 13080
rect 19544 13010 19554 13080
rect 19950 12900 20276 13192
rect 20594 12900 21008 13194
rect 21042 13018 21052 13076
rect 23024 13018 23034 13076
rect 19950 12898 23024 12900
rect 4770 12816 4780 12878
rect 6568 12816 6578 12878
rect 7996 12834 9172 12898
rect 11542 12834 11808 12898
rect 14178 12834 14188 12898
rect 17642 12896 21052 12898
rect 14526 12838 14536 12896
rect 16910 12838 17172 12896
rect 19546 12840 21052 12896
rect 23024 12840 23034 12898
rect 19546 12838 19556 12840
rect 4772 12754 4782 12756
rect 3772 12704 4782 12754
rect 3772 12518 4398 12704
rect 4772 12702 4782 12704
rect 6570 12702 6580 12756
rect 4768 12580 4778 12642
rect 6568 12580 6578 12642
rect 7996 12544 8448 12834
rect 9162 12654 9172 12724
rect 11540 12654 11550 12724
rect 11798 12654 11808 12724
rect 14176 12654 14186 12724
rect 14530 12654 14540 12724
rect 16908 12654 16918 12724
rect 17166 12654 17176 12724
rect 19544 12654 19554 12724
rect 4772 12518 4782 12520
rect 3772 12468 4782 12518
rect 3772 12282 4398 12468
rect 4772 12466 4782 12468
rect 6570 12466 6580 12520
rect 7996 12480 9172 12544
rect 11542 12480 11808 12544
rect 14178 12480 14188 12544
rect 19950 12542 20276 12840
rect 20594 12542 21008 12840
rect 21042 12662 21052 12720
rect 23024 12662 23034 12720
rect 14526 12482 14536 12540
rect 16910 12482 17172 12540
rect 19546 12538 19556 12540
rect 19950 12538 21052 12542
rect 19546 12484 21052 12538
rect 23024 12484 23034 12542
rect 19546 12482 23024 12484
rect 17594 12480 20276 12482
rect 4770 12344 4780 12406
rect 6568 12344 6578 12406
rect 4772 12282 4782 12284
rect 3772 12232 4782 12282
rect 3772 12044 4398 12232
rect 4772 12230 4782 12232
rect 6570 12230 6580 12284
rect 7996 12186 8448 12480
rect 9162 12298 9172 12368
rect 11540 12298 11550 12368
rect 11798 12298 11808 12368
rect 14176 12298 14186 12368
rect 14530 12298 14540 12368
rect 16908 12298 16918 12368
rect 17168 12298 17178 12368
rect 19546 12298 19556 12368
rect 19950 12188 20276 12480
rect 20594 12188 21008 12482
rect 21042 12306 21052 12364
rect 23024 12306 23034 12364
rect 19950 12186 23024 12188
rect 4770 12108 4780 12170
rect 6568 12108 6578 12170
rect 7996 12122 9172 12186
rect 11542 12122 11808 12186
rect 14178 12122 14188 12186
rect 19950 12184 21052 12186
rect 14526 12126 14536 12184
rect 16910 12126 17172 12184
rect 19546 12128 21052 12184
rect 23024 12128 23034 12186
rect 19546 12126 20276 12128
rect 4772 12044 4782 12048
rect 3772 11994 4782 12044
rect 6570 11994 6580 12048
rect 3772 11810 4398 11994
rect 4770 11872 4780 11934
rect 6568 11872 6578 11934
rect 7996 11830 8448 12122
rect 9162 11942 9172 12012
rect 11540 11942 11550 12012
rect 11798 11942 11808 12012
rect 14176 11942 14186 12012
rect 14530 11942 14540 12012
rect 16908 11942 16918 12012
rect 17168 11942 17178 12012
rect 19546 11942 19556 12012
rect 19950 11830 20276 12126
rect 20594 11830 21008 12128
rect 21042 11950 21052 12008
rect 23024 11950 23034 12008
rect 4772 11810 4782 11812
rect 3772 11760 4782 11810
rect 3772 11574 4398 11760
rect 4772 11758 4782 11760
rect 6570 11758 6580 11812
rect 7996 11766 9172 11830
rect 11542 11766 11808 11830
rect 14178 11766 14188 11830
rect 19950 11828 21052 11830
rect 14526 11770 14536 11828
rect 16910 11770 17172 11828
rect 19546 11772 21052 11828
rect 23024 11772 23034 11830
rect 19546 11770 23024 11772
rect 4768 11636 4778 11698
rect 6568 11636 6578 11698
rect 4772 11574 4782 11576
rect 3772 11524 4782 11574
rect 3772 11338 4398 11524
rect 4772 11522 4782 11524
rect 6570 11522 6580 11576
rect 7996 11476 8448 11766
rect 9160 11586 9170 11656
rect 11538 11586 11548 11656
rect 11798 11586 11808 11656
rect 14176 11586 14186 11656
rect 14530 11586 14540 11656
rect 16908 11586 16918 11656
rect 17166 11586 17176 11656
rect 19544 11586 19554 11656
rect 19950 11476 20276 11770
rect 20594 11476 21008 11770
rect 21042 11594 21052 11652
rect 23024 11594 23034 11652
rect 4768 11400 4778 11462
rect 6568 11400 6578 11462
rect 7996 11412 9172 11476
rect 11542 11412 11808 11476
rect 14178 11412 14188 11476
rect 19950 11474 23024 11476
rect 14526 11414 14536 11472
rect 16910 11414 17172 11472
rect 19546 11470 19556 11472
rect 19950 11470 21052 11474
rect 19546 11416 21052 11470
rect 23024 11416 23034 11474
rect 19546 11414 20276 11416
rect 17614 11412 20276 11414
rect 4772 11338 4782 11340
rect 3772 11288 4782 11338
rect 3772 11102 4398 11288
rect 4772 11286 4782 11288
rect 6570 11286 6580 11340
rect 4770 11164 4780 11226
rect 6568 11164 6578 11226
rect 7996 11120 8448 11412
rect 9160 11230 9170 11300
rect 11538 11230 11548 11300
rect 11798 11230 11808 11300
rect 14176 11230 14186 11300
rect 14530 11230 14540 11300
rect 16908 11230 16918 11300
rect 17166 11230 17176 11300
rect 19544 11230 19554 11300
rect 19950 11120 20276 11412
rect 20594 11120 21008 11416
rect 21042 11238 21052 11296
rect 23024 11238 23034 11296
rect 4772 11102 4782 11104
rect 3772 11052 4782 11102
rect 3772 10864 4398 11052
rect 4772 11050 4782 11052
rect 6570 11050 6580 11104
rect 7996 11056 9172 11120
rect 11542 11056 11808 11120
rect 14178 11056 14188 11120
rect 19950 11118 23024 11120
rect 19950 11116 21052 11118
rect 14526 11058 14536 11116
rect 16910 11058 17172 11116
rect 19546 11060 21052 11116
rect 23024 11060 23034 11118
rect 19546 11058 20276 11060
rect 4770 10928 4780 10990
rect 6568 10928 6578 10990
rect 4772 10864 4782 10868
rect 3772 10814 4782 10864
rect 6570 10814 6580 10868
rect 3772 10630 4398 10814
rect 7996 10764 8448 11056
rect 9160 10874 9170 10944
rect 11538 10874 11548 10944
rect 11798 10874 11808 10944
rect 14176 10874 14186 10944
rect 14530 10876 14540 10946
rect 16908 10876 16918 10946
rect 17166 10874 17176 10944
rect 19544 10874 19554 10944
rect 19950 10764 20276 11058
rect 20594 10764 21008 11060
rect 21042 10882 21052 10940
rect 23024 10882 23034 10940
rect 4770 10692 4780 10754
rect 6568 10692 6578 10754
rect 7996 10700 9172 10764
rect 11542 10700 11808 10764
rect 14178 10700 14188 10764
rect 19950 10762 23024 10764
rect 14526 10702 14536 10760
rect 16910 10702 17172 10760
rect 19546 10758 19556 10760
rect 19950 10758 21052 10762
rect 19546 10704 21052 10758
rect 23024 10704 23034 10762
rect 19546 10702 20276 10704
rect 17620 10700 20276 10702
rect 4772 10630 4782 10632
rect 3772 10580 4782 10630
rect 3772 10394 4398 10580
rect 4772 10578 4782 10580
rect 6570 10578 6580 10632
rect 4770 10456 4780 10518
rect 6568 10456 6578 10518
rect 7996 10408 8448 10700
rect 9160 10518 9170 10588
rect 11538 10518 11548 10588
rect 11798 10518 11808 10588
rect 14176 10518 14186 10588
rect 14528 10516 14538 10586
rect 16906 10516 16916 10586
rect 17166 10518 17176 10588
rect 19544 10518 19554 10588
rect 19950 10408 20276 10700
rect 20594 10408 21008 10704
rect 21042 10526 21052 10584
rect 23024 10526 23034 10584
rect 4772 10394 4782 10396
rect 3772 10344 4782 10394
rect 3772 10158 4398 10344
rect 4772 10342 4782 10344
rect 6570 10342 6580 10396
rect 7996 10344 9170 10408
rect 11540 10344 11808 10408
rect 14178 10344 14188 10408
rect 19950 10406 23024 10408
rect 17620 10404 21052 10406
rect 14526 10346 14536 10404
rect 16910 10346 17172 10404
rect 19546 10348 21052 10404
rect 23024 10348 23034 10406
rect 19546 10346 19556 10348
rect 4768 10220 4778 10282
rect 6568 10220 6578 10282
rect 4772 10158 4782 10160
rect 3772 10108 4782 10158
rect 3772 9922 4398 10108
rect 4772 10106 4782 10108
rect 6570 10106 6580 10160
rect 7996 10052 8448 10344
rect 9160 10160 9170 10232
rect 11538 10160 11548 10232
rect 11798 10162 11808 10232
rect 14176 10162 14186 10232
rect 14530 10162 14540 10232
rect 16908 10162 16918 10232
rect 17166 10162 17176 10232
rect 19544 10162 19554 10232
rect 4768 9984 4778 10046
rect 6568 9984 6578 10046
rect 7996 9988 9172 10052
rect 11542 9988 11808 10052
rect 14178 9988 14188 10052
rect 19950 10050 20276 10348
rect 20594 10050 21008 10348
rect 21042 10170 21052 10228
rect 23024 10170 23034 10228
rect 19950 10048 21052 10050
rect 14526 9990 14536 10048
rect 16910 9990 17172 10048
rect 19546 9992 21052 10048
rect 23024 9992 23034 10050
rect 19546 9990 23024 9992
rect 4772 9922 4782 9924
rect 3772 9872 4782 9922
rect 3772 9686 4398 9872
rect 4772 9870 4782 9872
rect 6570 9870 6580 9924
rect 4770 9748 4780 9810
rect 6568 9748 6578 9810
rect 7996 9696 8448 9988
rect 9160 9806 9170 9876
rect 11538 9806 11548 9876
rect 11798 9806 11808 9876
rect 14176 9806 14186 9876
rect 14530 9806 14540 9876
rect 16908 9806 16918 9876
rect 17166 9806 17176 9876
rect 19544 9806 19554 9876
rect 4772 9686 4782 9688
rect 3772 9636 4782 9686
rect 3772 9450 4398 9636
rect 4772 9634 4782 9636
rect 6570 9634 6580 9688
rect 7996 9632 9172 9696
rect 11542 9632 11808 9696
rect 14178 9632 14188 9696
rect 19950 9694 20276 9990
rect 20594 9694 21008 9990
rect 21042 9814 21052 9872
rect 23024 9814 23034 9872
rect 19950 9692 21052 9694
rect 14526 9634 14536 9692
rect 16910 9634 17172 9692
rect 19546 9636 21052 9692
rect 23024 9636 23034 9694
rect 19546 9634 23024 9636
rect 4768 9512 4778 9574
rect 6568 9512 6578 9574
rect 4772 9450 4782 9452
rect 3772 9400 4782 9450
rect 3772 9214 4398 9400
rect 4772 9398 4782 9400
rect 6570 9398 6580 9452
rect 7996 9340 8448 9632
rect 9162 9450 9172 9520
rect 11540 9450 11550 9520
rect 11798 9450 11808 9520
rect 14176 9450 14186 9520
rect 14528 9450 14538 9520
rect 16906 9450 16916 9520
rect 17166 9450 17176 9520
rect 19544 9450 19554 9520
rect 9162 9340 9172 9342
rect 4770 9276 4780 9338
rect 6568 9276 6578 9338
rect 7996 9278 9172 9340
rect 11542 9340 11552 9342
rect 11542 9278 11808 9340
rect 7996 9276 11808 9278
rect 14178 9276 14188 9340
rect 19950 9338 20276 9634
rect 20594 9338 21008 9634
rect 21042 9458 21052 9516
rect 23024 9458 23034 9516
rect 14526 9280 14536 9338
rect 16910 9336 16920 9338
rect 16910 9280 17172 9336
rect 14538 9278 17172 9280
rect 19546 9334 19556 9336
rect 19950 9334 21052 9338
rect 19546 9280 21052 9334
rect 23024 9280 23034 9338
rect 19546 9278 23024 9280
rect 17618 9276 20276 9278
rect 4770 9214 4780 9216
rect 3772 9164 4780 9214
rect 3772 8976 4398 9164
rect 4770 9162 4780 9164
rect 6568 9162 6578 9216
rect 4770 9100 4780 9102
rect 4768 9038 4778 9100
rect 6568 9038 6578 9102
rect 7996 8982 8448 9276
rect 9162 9094 9172 9164
rect 11540 9094 11550 9164
rect 11800 9094 11810 9164
rect 14178 9094 14188 9164
rect 14528 9094 14538 9164
rect 16906 9094 16916 9164
rect 17166 9094 17176 9164
rect 19544 9094 19554 9164
rect 19950 8982 20276 9276
rect 20594 8982 21008 9278
rect 21042 9102 21052 9160
rect 23024 9102 23034 9160
rect 4770 8976 4780 8980
rect 3772 8926 4780 8976
rect 6568 8926 6578 8980
rect 3772 8742 4398 8926
rect 7996 8918 9172 8982
rect 11542 8918 11808 8982
rect 14178 8918 14188 8982
rect 14526 8922 14536 8980
rect 16910 8922 17172 8980
rect 19546 8978 19556 8980
rect 19950 8978 21052 8982
rect 19546 8924 21052 8978
rect 23024 8924 23034 8982
rect 19546 8922 23024 8924
rect 17616 8920 20276 8922
rect 4770 8866 4780 8868
rect 4768 8804 4778 8866
rect 6568 8804 6578 8868
rect 4770 8742 4780 8744
rect 3772 8692 4780 8742
rect 3772 8280 4398 8692
rect 4770 8690 4780 8692
rect 6568 8690 6578 8744
rect 4770 8568 4780 8632
rect 6568 8568 6578 8632
rect 7996 8628 8448 8918
rect 9162 8736 9172 8806
rect 11540 8736 11550 8806
rect 11800 8738 11810 8808
rect 14178 8738 14188 8808
rect 14528 8736 14538 8806
rect 16906 8736 16916 8806
rect 17166 8738 17176 8808
rect 19544 8738 19554 8808
rect 19950 8628 20276 8920
rect 20594 8628 21008 8922
rect 21042 8746 21052 8804
rect 23024 8746 23034 8804
rect 7996 8626 11808 8628
rect 7996 8564 9172 8626
rect 4778 8280 4788 8282
rect 3772 8230 4788 8280
rect 3772 8042 4398 8230
rect 4778 8224 4788 8230
rect 6568 8224 6578 8282
rect 7996 8272 8448 8564
rect 9162 8562 9172 8564
rect 11542 8564 11808 8626
rect 14178 8564 14188 8628
rect 19950 8626 23024 8628
rect 19950 8624 21052 8626
rect 14524 8566 14534 8624
rect 16908 8566 17172 8624
rect 19546 8568 21052 8624
rect 23024 8568 23034 8626
rect 19546 8566 20276 8568
rect 11542 8562 11552 8564
rect 9162 8382 9172 8452
rect 11540 8382 11550 8452
rect 11798 8382 11808 8452
rect 14176 8382 14186 8452
rect 14528 8382 14538 8452
rect 16906 8382 16916 8452
rect 17166 8382 17176 8452
rect 19544 8382 19554 8452
rect 7996 8208 9172 8272
rect 11542 8208 11806 8272
rect 14176 8208 14186 8272
rect 19950 8270 20276 8566
rect 20594 8270 21008 8568
rect 21044 8390 21054 8448
rect 23026 8390 23036 8448
rect 19950 8268 21052 8270
rect 14526 8210 14536 8268
rect 16910 8210 17172 8268
rect 19546 8212 21052 8268
rect 23024 8212 23034 8270
rect 19546 8210 23024 8212
rect 4778 8042 4788 8046
rect 3772 7992 4788 8042
rect 3772 7808 4398 7992
rect 4778 7988 4788 7992
rect 6568 7988 6578 8046
rect 7996 7916 8448 8208
rect 9162 8026 9172 8096
rect 11540 8026 11550 8096
rect 11800 8026 11810 8096
rect 14178 8026 14188 8096
rect 14530 8026 14540 8096
rect 16908 8026 16918 8096
rect 17166 8026 17176 8096
rect 19544 8026 19554 8096
rect 7996 7852 9172 7916
rect 11542 7914 14178 7916
rect 19950 7914 20276 8210
rect 20594 7914 21008 8210
rect 21042 8034 21052 8092
rect 23024 8034 23034 8092
rect 11542 7852 11808 7914
rect 4778 7808 4788 7810
rect 3772 7758 4788 7808
rect 3772 7640 4398 7758
rect 4778 7752 4788 7758
rect 6568 7752 6578 7810
rect 3772 7638 4394 7640
rect 3772 3110 4380 7638
rect 220 2496 580 2506
rect 1996 2184 4380 3110
rect 7996 7560 8448 7852
rect 11798 7850 11808 7852
rect 14178 7850 14188 7914
rect 14526 7854 14536 7912
rect 16910 7854 17172 7912
rect 19546 7910 19556 7912
rect 19950 7910 21052 7914
rect 19546 7856 21052 7910
rect 23024 7856 23034 7914
rect 19546 7854 23024 7856
rect 17628 7852 20276 7854
rect 9162 7670 9172 7740
rect 11540 7670 11550 7740
rect 11798 7670 11808 7740
rect 14176 7670 14186 7740
rect 14530 7672 14540 7742
rect 16908 7672 16918 7742
rect 17166 7670 17176 7740
rect 19544 7670 19554 7740
rect 19950 7560 20276 7852
rect 20594 7560 21008 7854
rect 21042 7678 21052 7736
rect 23024 7678 23034 7736
rect 7996 7496 9172 7560
rect 11542 7496 11808 7560
rect 14178 7496 14188 7560
rect 19950 7558 23024 7560
rect 17638 7556 21052 7558
rect 14526 7498 14536 7556
rect 16910 7498 17172 7556
rect 19546 7500 21052 7556
rect 23024 7500 23034 7558
rect 19546 7498 19556 7500
rect 7996 7204 8448 7496
rect 9162 7314 9172 7384
rect 11540 7314 11550 7384
rect 11798 7314 11808 7384
rect 14176 7314 14186 7384
rect 14530 7314 14540 7384
rect 16908 7314 16918 7384
rect 17166 7314 17176 7384
rect 19544 7314 19554 7384
rect 7996 7140 9172 7204
rect 11542 7140 11808 7204
rect 14178 7140 14188 7204
rect 19950 7202 20276 7500
rect 20594 7202 21008 7500
rect 21042 7322 21052 7380
rect 23024 7322 23034 7380
rect 19950 7200 21052 7202
rect 14526 7142 14536 7200
rect 16910 7198 21052 7200
rect 16910 7142 17172 7198
rect 17162 7140 17172 7142
rect 19546 7144 21052 7198
rect 23024 7144 23034 7202
rect 19546 7142 23024 7144
rect 19546 7140 19556 7142
rect 7996 6848 8448 7140
rect 9162 6958 9172 7028
rect 11540 6958 11550 7028
rect 11800 6958 11810 7028
rect 14178 6958 14188 7028
rect 14530 6956 14540 7026
rect 16908 6956 16918 7026
rect 17166 6958 17176 7028
rect 19544 6958 19554 7028
rect 19950 6848 20276 7142
rect 20594 6848 21008 7142
rect 21042 6966 21052 7024
rect 23024 6966 23034 7024
rect 7996 6784 9172 6848
rect 11542 6784 11808 6848
rect 14178 6784 14188 6848
rect 19950 6846 21052 6848
rect 17628 6844 21052 6846
rect 14526 6786 14536 6844
rect 16910 6786 17172 6844
rect 19546 6790 21052 6844
rect 23024 6790 23034 6848
rect 19546 6788 23024 6790
rect 19546 6786 19556 6788
rect 7996 6492 8448 6784
rect 9162 6602 9172 6672
rect 11540 6602 11550 6672
rect 11798 6602 11808 6672
rect 14176 6602 14186 6672
rect 14530 6602 14540 6672
rect 16908 6602 16918 6672
rect 17166 6602 17176 6672
rect 19544 6602 19554 6672
rect 7996 6428 9172 6492
rect 11542 6490 14178 6492
rect 19950 6490 20276 6788
rect 20594 6490 21008 6788
rect 21042 6610 21052 6668
rect 23024 6610 23034 6668
rect 11542 6428 11808 6490
rect 7996 6136 8448 6428
rect 11798 6426 11808 6428
rect 14178 6426 14188 6490
rect 19950 6488 21052 6490
rect 14526 6430 14536 6488
rect 16910 6430 17172 6488
rect 19546 6432 21052 6488
rect 23024 6432 23034 6490
rect 19546 6430 23024 6432
rect 9162 6246 9172 6316
rect 11540 6246 11550 6316
rect 11800 6246 11810 6316
rect 14178 6246 14188 6316
rect 14530 6246 14540 6316
rect 16908 6246 16918 6316
rect 17166 6246 17176 6316
rect 19544 6246 19554 6316
rect 19950 6136 20276 6430
rect 20594 6136 21008 6430
rect 21042 6254 21052 6312
rect 23024 6254 23034 6312
rect 7996 6072 9172 6136
rect 11542 6072 11808 6136
rect 14178 6072 14188 6136
rect 19950 6134 23024 6136
rect 19950 6132 21052 6134
rect 14526 6074 14536 6132
rect 16910 6074 17172 6132
rect 19546 6076 21052 6132
rect 23024 6076 23034 6134
rect 19546 6074 20276 6076
rect 7996 5778 8448 6072
rect 9160 5890 9170 5960
rect 11538 5890 11548 5960
rect 11800 5890 11810 5960
rect 14178 5890 14188 5960
rect 14530 5892 14540 5962
rect 16908 5892 16918 5962
rect 17166 5890 17176 5960
rect 19544 5890 19554 5960
rect 19950 5780 20276 6074
rect 20594 5780 21008 6076
rect 21042 5898 21052 5956
rect 23024 5898 23034 5956
rect 19950 5778 23024 5780
rect 7996 5714 9172 5778
rect 11542 5714 11808 5778
rect 14178 5714 14188 5778
rect 19950 5776 21052 5778
rect 14526 5718 14536 5776
rect 16910 5718 17172 5776
rect 19546 5720 21052 5776
rect 23024 5720 23034 5778
rect 19546 5718 20276 5720
rect 7996 5422 8448 5714
rect 9162 5534 9172 5604
rect 11540 5534 11550 5604
rect 11798 5534 11808 5604
rect 14176 5534 14186 5604
rect 14530 5534 14540 5604
rect 16908 5534 16918 5604
rect 17166 5534 17176 5604
rect 19544 5534 19554 5604
rect 19950 5424 20276 5718
rect 20594 5424 21008 5720
rect 21042 5542 21052 5600
rect 23024 5542 23034 5600
rect 19950 5422 23024 5424
rect 7996 5358 9172 5422
rect 11542 5358 11808 5422
rect 14178 5358 14188 5422
rect 19950 5420 21052 5422
rect 14526 5362 14536 5420
rect 16910 5362 17172 5420
rect 19546 5364 21052 5420
rect 23024 5364 23034 5422
rect 19546 5362 20276 5364
rect 7996 5066 8448 5358
rect 9162 5176 9172 5246
rect 11540 5176 11550 5246
rect 11798 5178 11808 5248
rect 14176 5178 14186 5248
rect 14530 5176 14540 5246
rect 16908 5176 16918 5246
rect 17166 5178 17176 5248
rect 19544 5178 19554 5248
rect 19950 5068 20276 5362
rect 20594 5068 21008 5364
rect 21042 5186 21052 5244
rect 23024 5186 23034 5244
rect 7996 5002 9172 5066
rect 11542 5002 11806 5066
rect 14176 5002 14186 5066
rect 19950 5064 21052 5068
rect 14526 5006 14536 5064
rect 16910 5006 17172 5064
rect 19546 5010 21052 5064
rect 23024 5010 23034 5068
rect 19546 5008 23024 5010
rect 19546 5006 20276 5008
rect 7996 4712 8448 5002
rect 9162 4822 9172 4892
rect 11542 4822 11552 4892
rect 11798 4822 11808 4892
rect 14176 4822 14186 4892
rect 14530 4822 14540 4892
rect 16908 4822 16918 4892
rect 17166 4822 17176 4892
rect 19544 4822 19554 4892
rect 7996 4648 9172 4712
rect 11542 4648 11806 4712
rect 14176 4648 14186 4712
rect 19950 4710 20276 5006
rect 20594 4710 21008 5008
rect 21042 4830 21052 4888
rect 23024 4830 23034 4888
rect 19950 4708 21052 4710
rect 14526 4650 14536 4708
rect 16910 4650 17172 4708
rect 19546 4652 21052 4708
rect 23024 4652 23034 4710
rect 19546 4650 23024 4652
rect 7996 4356 8448 4648
rect 9162 4466 9172 4536
rect 11540 4466 11550 4536
rect 11798 4466 11808 4536
rect 14176 4466 14186 4536
rect 14530 4466 14540 4536
rect 16908 4466 16918 4536
rect 17166 4466 17176 4536
rect 19544 4466 19554 4536
rect 19950 4356 20276 4650
rect 20594 4356 21008 4650
rect 21042 4474 21052 4532
rect 23024 4474 23034 4532
rect 7996 4292 9172 4356
rect 11542 4354 14178 4356
rect 19950 4354 23024 4356
rect 11542 4292 11808 4354
rect 7996 3998 8448 4292
rect 11798 4290 11808 4292
rect 14178 4290 14188 4354
rect 19950 4352 21052 4354
rect 14526 4294 14536 4352
rect 16910 4294 17172 4352
rect 19546 4296 21052 4352
rect 23024 4296 23034 4354
rect 19546 4294 20276 4296
rect 9162 4110 9172 4180
rect 11540 4110 11550 4180
rect 11798 4110 11808 4180
rect 14176 4110 14186 4180
rect 14530 4110 14540 4180
rect 16908 4110 16918 4180
rect 17166 4110 17176 4180
rect 19544 4110 19554 4180
rect 19950 4000 20276 4294
rect 20594 4000 21008 4296
rect 21042 4118 21052 4176
rect 23024 4118 23034 4176
rect 7996 3934 9172 3998
rect 11542 3934 11808 3998
rect 14178 3934 14188 3998
rect 19950 3996 21052 4000
rect 14526 3938 14536 3996
rect 16910 3994 21052 3996
rect 16910 3938 17172 3994
rect 17162 3936 17172 3938
rect 19546 3942 21052 3994
rect 23024 3942 23034 4000
rect 19546 3940 23024 3942
rect 19546 3938 20276 3940
rect 19546 3936 19556 3938
rect 7996 3642 8448 3934
rect 9162 3754 9172 3824
rect 11540 3754 11550 3824
rect 11798 3754 11808 3824
rect 14176 3754 14186 3824
rect 14530 3754 14540 3824
rect 16908 3754 16918 3824
rect 17166 3754 17176 3824
rect 19544 3754 19554 3824
rect 7996 3578 9172 3642
rect 11542 3578 11806 3642
rect 14176 3578 14186 3642
rect 19950 3640 20276 3938
rect 20594 3640 21008 3940
rect 21042 3762 21052 3820
rect 23024 3762 23034 3820
rect 21042 3640 21052 3642
rect 14526 3582 14536 3640
rect 16910 3582 17172 3640
rect 19546 3584 21052 3640
rect 23024 3584 23034 3642
rect 19546 3582 23024 3584
rect 19950 3580 23024 3582
rect 7996 3288 8448 3578
rect 9162 3398 9172 3468
rect 11540 3398 11550 3468
rect 11798 3398 11808 3468
rect 14176 3398 14186 3468
rect 14530 3396 14540 3466
rect 16908 3396 16918 3466
rect 17166 3398 17176 3468
rect 19544 3398 19554 3468
rect 19950 3288 20276 3580
rect 20594 3288 21008 3580
rect 21042 3406 21052 3464
rect 23024 3406 23034 3464
rect 7996 3224 9172 3288
rect 11542 3224 11808 3288
rect 14178 3224 14188 3288
rect 19950 3286 23024 3288
rect 19950 3284 21052 3286
rect 14526 3226 14536 3284
rect 16910 3226 17170 3284
rect 19544 3228 21052 3284
rect 23024 3228 23034 3286
rect 19544 3226 20276 3228
rect 7996 2932 8448 3224
rect 9162 3042 9172 3112
rect 11540 3042 11550 3112
rect 11798 3042 11808 3112
rect 14176 3042 14186 3112
rect 14530 3042 14540 3112
rect 16908 3042 16918 3112
rect 17166 3042 17176 3112
rect 19544 3042 19554 3112
rect 7996 2868 9172 2932
rect 11542 2868 11806 2932
rect 14176 2868 14186 2932
rect 19950 2930 20276 3226
rect 20594 2930 21008 3228
rect 21042 3050 21052 3108
rect 23024 3050 23034 3108
rect 19950 2928 21052 2930
rect 14526 2870 14536 2928
rect 16910 2870 17170 2928
rect 19544 2872 21052 2928
rect 23024 2872 23034 2930
rect 19544 2870 23024 2872
rect 7996 2774 8448 2868
rect 19950 2762 20276 2870
rect 20594 2842 21008 2870
rect 20594 2840 20858 2842
rect 23241 2734 25116 27192
rect 25640 2734 27492 40588
rect 11182 2286 12192 2296
rect 580 1296 4380 2184
rect 220 1038 580 1048
rect 1996 1000 4380 1296
rect 6242 2272 7252 2282
rect 11182 1284 12192 1294
rect 16524 2286 17534 2296
rect 23241 1960 27492 2734
rect 16524 1284 17534 1294
rect 6242 1270 7252 1280
rect 23242 1000 27492 1960
<< via2 >>
rect 23738 43240 27086 43860
rect 20656 40396 23026 40460
rect 20656 40160 23026 40224
rect 20654 39924 23024 39988
rect 20654 39688 23024 39752
rect 20656 39452 23026 39516
rect 20654 39214 23024 39278
rect 20656 38978 23026 39042
rect 20654 38746 23024 38810
rect 20656 38506 23026 38570
rect 20654 38270 23024 38334
rect 3018 38138 4792 38204
rect 20654 38034 23024 38098
rect 3018 37902 4792 37968
rect 20656 37798 23026 37862
rect 3018 37666 4792 37732
rect 20656 37562 23026 37626
rect 3018 37430 4792 37496
rect 20656 37326 23026 37390
rect 3018 37194 4792 37260
rect 20654 37092 23024 37156
rect 3018 36958 4792 37024
rect 20658 36856 23028 36920
rect 3018 36722 4792 36788
rect 20656 36618 23026 36682
rect 3018 36486 4792 36552
rect 20658 36382 23028 36446
rect 3018 36250 4792 36316
rect 20658 36146 23028 36210
rect 3018 36014 4792 36080
rect 20658 35912 23028 35976
rect 3018 35778 4792 35844
rect 20654 35674 23024 35738
rect 3018 35542 4792 35608
rect 20654 35436 23024 35500
rect 3018 35306 4792 35372
rect 20656 35202 23026 35266
rect 3018 35070 4792 35136
rect 20656 34966 23026 35030
rect 3018 34834 4792 34900
rect 20658 34730 23028 34794
rect 3018 34598 4792 34664
rect 20654 34496 23024 34560
rect 3018 34362 4792 34428
rect 20654 34258 23024 34322
rect 3018 34126 4792 34192
rect 20656 34024 23026 34088
rect 3018 33890 4792 33956
rect 20656 33786 23026 33850
rect 3018 33654 4792 33720
rect 20656 33550 23026 33614
rect 3018 33418 4792 33484
rect 20656 33316 23026 33380
rect 3018 33182 4792 33248
rect 20656 33080 23026 33144
rect 3018 32946 4792 33012
rect 20656 32842 23026 32906
rect 3018 32710 4792 32776
rect 20658 32608 23028 32672
rect 3018 32474 4792 32540
rect 20658 32374 23028 32438
rect 3018 32238 4792 32304
rect 20656 32134 23026 32198
rect 3018 32002 4792 32068
rect 20656 31900 23026 31964
rect 3016 31766 4790 31832
rect 20656 31662 23026 31726
rect 3018 31530 4792 31596
rect 20656 31428 23026 31492
rect 3018 31294 4792 31360
rect 20656 31192 23026 31256
rect 3018 31060 4792 31120
rect 20654 30956 23024 31020
rect 20656 30718 23026 30782
rect 20656 30482 23026 30546
rect 20656 30248 23026 30312
rect 20656 30010 23026 30074
rect 20658 29776 23028 29840
rect 18478 22294 18982 22684
rect 19814 22660 19974 22772
rect 19810 21030 19970 21144
rect 9172 20486 9174 20556
rect 9174 20486 11540 20556
rect 11808 20486 14176 20556
rect 14540 20488 16908 20558
rect 17176 20486 19544 20556
rect 9172 20130 11540 20200
rect 11808 20130 14176 20200
rect 14540 20130 16908 20200
rect 17176 20130 19544 20200
rect 9172 19774 11540 19844
rect 11808 19774 14176 19844
rect 14540 19774 16908 19844
rect 17176 19774 19544 19844
rect 9172 19420 11540 19490
rect 11808 19418 14176 19488
rect 14540 19416 16908 19486
rect 17176 19416 19544 19486
rect 9172 19062 11540 19132
rect 11808 19062 14176 19132
rect 14540 19062 16908 19132
rect 17176 19062 19544 19132
rect 9172 18706 11540 18776
rect 11808 18706 14176 18776
rect 14540 18706 16908 18776
rect 17176 18706 19544 18776
rect 9172 18350 11540 18420
rect 11808 18350 14176 18420
rect 14540 18350 16908 18420
rect 17176 18350 19544 18420
rect 9172 17994 11540 18064
rect 11808 17994 14176 18064
rect 14540 17994 16908 18064
rect 17176 17994 19544 18064
rect 9172 17638 11540 17708
rect 11808 17638 14176 17708
rect 14540 17638 16908 17708
rect 17176 17636 19544 17706
rect 9172 17350 11540 17352
rect 9172 17282 11540 17350
rect 11808 17282 14176 17352
rect 14540 17282 16908 17352
rect 17176 17282 19544 17352
rect 9172 16926 11540 16996
rect 11808 16926 14176 16996
rect 14540 16926 16908 16996
rect 17176 16926 19544 16996
rect 9172 16570 11540 16640
rect 11808 16570 14176 16640
rect 14540 16570 16908 16640
rect 17176 16570 19544 16640
rect 9172 16216 11540 16284
rect 9172 16214 11540 16216
rect 11808 16216 14176 16286
rect 14540 16214 16908 16284
rect 17176 16214 19544 16284
rect 9172 15858 11540 15928
rect 11808 15858 14176 15928
rect 14540 15856 16908 15926
rect 17176 15858 19544 15928
rect 4780 15648 6568 15710
rect 4780 15412 6568 15474
rect 9172 15502 11540 15572
rect 11808 15502 14176 15572
rect 14540 15502 16908 15572
rect 17176 15502 19544 15572
rect 4780 15176 6568 15238
rect 9172 15146 11540 15216
rect 11808 15146 14176 15216
rect 14540 15146 16908 15216
rect 17176 15146 19544 15216
rect 4780 14940 6568 15002
rect 4780 14704 6568 14766
rect 9172 14790 11540 14860
rect 11808 14790 14176 14860
rect 14540 14790 16908 14860
rect 17176 14790 19544 14860
rect 4780 14468 6568 14530
rect 9172 14434 11540 14504
rect 11808 14434 14176 14504
rect 14540 14434 16908 14504
rect 17176 14434 19544 14504
rect 4780 14232 6568 14294
rect 4780 13996 6566 14058
rect 6566 13996 6568 14058
rect 9172 14078 11540 14148
rect 11808 14078 14176 14148
rect 14540 14076 16908 14146
rect 17176 14078 19544 14148
rect 21054 24992 23024 25056
rect 21054 24636 23024 24700
rect 21054 24278 23024 24342
rect 21054 23922 23024 23986
rect 21052 23568 23022 23632
rect 21054 23210 23024 23274
rect 21054 22856 23024 22920
rect 21054 22498 23024 22562
rect 21054 22142 23024 22206
rect 21054 21788 23024 21852
rect 21054 21430 23024 21494
rect 21054 21076 23024 21140
rect 21052 20718 23022 20782
rect 21054 20360 23024 20424
rect 21052 20008 23022 20072
rect 21054 19650 23024 19714
rect 21052 19296 23022 19360
rect 21054 18938 23024 19002
rect 21052 18582 23022 18646
rect 21054 18226 23024 18290
rect 21054 17870 23024 17934
rect 21054 17514 23024 17578
rect 21054 17158 23024 17222
rect 21054 16802 23024 16866
rect 21052 16446 23022 16510
rect 21054 16090 23024 16154
rect 21054 15736 23024 15800
rect 21054 15378 23024 15442
rect 21054 15022 23024 15086
rect 21054 14668 23024 14732
rect 21054 14310 23024 14374
rect 4780 13760 6568 13822
rect 9172 13722 11540 13792
rect 11808 13722 14176 13792
rect 14540 13722 16908 13792
rect 17176 13722 19544 13792
rect 4780 13524 6568 13586
rect 21052 13730 23024 13788
rect 4780 13288 6568 13350
rect 9172 13366 11540 13436
rect 11808 13366 14176 13436
rect 14540 13366 16908 13436
rect 17176 13366 19544 13436
rect 21052 13374 23024 13432
rect 4780 13052 6568 13114
rect 9172 13010 11540 13080
rect 11808 13010 14176 13080
rect 14540 13010 16908 13080
rect 17176 13010 19544 13080
rect 21052 13018 23024 13076
rect 4780 12816 6568 12878
rect 4780 12580 6566 12642
rect 6566 12580 6568 12642
rect 9172 12654 11540 12724
rect 11808 12654 14176 12724
rect 14540 12654 16908 12724
rect 17176 12654 19544 12724
rect 21052 12662 23024 12720
rect 4780 12344 6568 12406
rect 9172 12298 11540 12368
rect 11808 12298 14176 12368
rect 14540 12298 16908 12368
rect 17178 12298 19546 12368
rect 21052 12306 23024 12364
rect 4780 12108 6568 12170
rect 4780 11872 6568 11934
rect 9172 11942 11540 12012
rect 11808 11942 14176 12012
rect 14540 11942 16908 12012
rect 17178 11942 19546 12012
rect 21052 11950 23024 12008
rect 4780 11636 6566 11698
rect 6566 11636 6568 11698
rect 9170 11586 11538 11656
rect 11808 11586 14176 11656
rect 14540 11586 16908 11656
rect 17176 11586 19544 11656
rect 21052 11594 23024 11652
rect 4780 11400 6566 11462
rect 6566 11400 6568 11462
rect 4780 11164 6568 11226
rect 9170 11230 11538 11300
rect 11808 11230 14176 11300
rect 14540 11230 16908 11300
rect 17176 11230 19544 11300
rect 21052 11238 23024 11296
rect 4780 10928 6568 10990
rect 9170 10874 11538 10944
rect 11808 10874 14176 10944
rect 14540 10876 16908 10946
rect 17176 10874 19544 10944
rect 21052 10882 23024 10940
rect 4780 10692 6568 10754
rect 4780 10456 6568 10518
rect 9170 10518 11538 10588
rect 11808 10518 14176 10588
rect 14538 10516 16906 10586
rect 17176 10518 19544 10588
rect 21052 10526 23024 10584
rect 4780 10220 6566 10282
rect 6566 10220 6568 10282
rect 9170 10230 11538 10232
rect 9170 10162 11538 10230
rect 11808 10162 14176 10232
rect 14540 10162 16908 10232
rect 17176 10162 19544 10232
rect 4780 9984 6566 10046
rect 6566 9984 6568 10046
rect 21052 10170 23024 10228
rect 4780 9748 6568 9810
rect 9170 9806 11538 9876
rect 11808 9806 14176 9876
rect 14540 9806 16908 9876
rect 17176 9806 19544 9876
rect 21052 9814 23024 9872
rect 4780 9512 6566 9574
rect 6566 9512 6568 9574
rect 9172 9450 11540 9520
rect 11808 9450 14176 9520
rect 14538 9450 16906 9520
rect 17176 9450 19544 9520
rect 4780 9276 6568 9338
rect 21052 9458 23024 9516
rect 4780 9100 6568 9102
rect 4780 9038 6566 9100
rect 6566 9038 6568 9100
rect 9172 9094 11540 9164
rect 11810 9094 14178 9164
rect 14538 9094 16906 9164
rect 17176 9094 19544 9164
rect 21052 9102 23024 9160
rect 4780 8866 6568 8868
rect 4780 8804 6566 8866
rect 6566 8804 6568 8866
rect 4780 8630 6568 8632
rect 4780 8568 6568 8630
rect 9172 8736 11540 8806
rect 11810 8738 14178 8808
rect 14538 8736 16906 8806
rect 17176 8738 19544 8808
rect 21052 8746 23024 8804
rect 9172 8382 11540 8452
rect 11808 8382 14176 8452
rect 14538 8382 16906 8452
rect 17176 8382 19544 8452
rect 21054 8390 23026 8448
rect 9172 8026 11540 8096
rect 11810 8026 14178 8096
rect 14540 8026 16908 8096
rect 17176 8026 19544 8096
rect 21052 8034 23024 8092
rect 220 1048 580 2496
rect 9172 7670 11540 7740
rect 11808 7670 14176 7740
rect 14540 7672 16908 7742
rect 17176 7670 19544 7740
rect 21052 7678 23024 7736
rect 9172 7314 11540 7384
rect 11808 7314 14176 7384
rect 14540 7314 16908 7384
rect 17176 7314 19544 7384
rect 21052 7322 23024 7380
rect 9172 6958 11540 7028
rect 11810 6958 14178 7028
rect 14540 6956 16908 7026
rect 17176 6958 19544 7028
rect 21052 6966 23024 7024
rect 9172 6602 11540 6672
rect 11808 6602 14176 6672
rect 14540 6602 16908 6672
rect 17176 6602 19544 6672
rect 21052 6610 23024 6668
rect 9172 6246 11540 6316
rect 11810 6246 14178 6316
rect 14540 6246 16908 6316
rect 17176 6246 19544 6316
rect 21052 6254 23024 6312
rect 9170 5890 11538 5960
rect 11810 5890 14178 5960
rect 14540 5892 16908 5962
rect 17176 5890 19544 5960
rect 21052 5898 23024 5956
rect 9172 5534 11540 5604
rect 11808 5534 14176 5604
rect 14540 5534 16908 5604
rect 17176 5534 19544 5604
rect 21052 5542 23024 5600
rect 9172 5176 11540 5246
rect 11808 5178 14176 5248
rect 14540 5176 16908 5246
rect 17176 5178 19544 5248
rect 21052 5186 23024 5244
rect 9172 4822 9174 4892
rect 9174 4822 11540 4892
rect 11808 4822 14176 4892
rect 14540 4822 16908 4892
rect 17176 4822 19544 4892
rect 21052 4830 23024 4888
rect 9172 4466 11540 4536
rect 11808 4466 14176 4536
rect 14540 4466 16908 4536
rect 17176 4466 19544 4536
rect 21052 4474 23024 4532
rect 9172 4110 11540 4180
rect 11808 4110 14176 4180
rect 14540 4110 16908 4180
rect 17176 4110 19544 4180
rect 21052 4118 23024 4176
rect 9172 3754 11540 3824
rect 11808 3754 14176 3824
rect 14540 3754 16908 3824
rect 17176 3754 19544 3824
rect 21052 3762 23024 3820
rect 9172 3398 11540 3468
rect 11808 3398 14176 3468
rect 14540 3396 16908 3466
rect 17176 3398 19544 3468
rect 21052 3406 23024 3464
rect 9172 3042 11540 3112
rect 11808 3042 14176 3112
rect 14540 3042 16908 3112
rect 17176 3042 19544 3112
rect 21052 3050 23024 3108
rect 25116 2734 25640 40588
rect 6242 1280 7252 2272
rect 11182 1294 12192 2286
rect 16524 1294 17534 2286
<< metal3 >>
rect 23260 43860 27492 44454
rect 3013 38204 4797 38214
rect 3013 38138 3018 38204
rect 4792 38202 4797 38204
rect 5224 38202 5754 38296
rect 4792 38168 5754 38202
rect 4792 38138 5342 38168
rect 3013 38136 5342 38138
rect 3013 38128 4797 38136
rect 3013 37970 4797 37978
rect 5224 37970 5342 38136
rect 3013 37968 5342 37970
rect 3013 37902 3018 37968
rect 4792 37904 5342 37968
rect 4792 37902 4797 37904
rect 3013 37892 4797 37902
rect 3013 37732 4797 37742
rect 5224 37732 5342 37904
rect 3013 37666 3018 37732
rect 4792 37666 5342 37732
rect 3013 37656 4797 37666
rect 3013 37498 4797 37506
rect 5224 37498 5342 37666
rect 3013 37496 5342 37498
rect 3013 37430 3018 37496
rect 4792 37432 5342 37496
rect 4792 37430 4797 37432
rect 3013 37420 4797 37430
rect 3013 37260 4797 37270
rect 5224 37260 5342 37432
rect 3013 37194 3018 37260
rect 4792 37194 5342 37260
rect 3013 37184 4797 37194
rect 3013 37024 4797 37034
rect 5224 37024 5342 37194
rect 3013 36958 3018 37024
rect 4792 36958 5342 37024
rect 3013 36948 4797 36958
rect 3013 36790 4797 36798
rect 5224 36790 5342 36958
rect 3013 36788 5342 36790
rect 3013 36722 3018 36788
rect 4792 36724 5342 36788
rect 4792 36722 4797 36724
rect 3013 36712 4797 36722
rect 3013 36552 4797 36562
rect 3013 36486 3018 36552
rect 4792 36550 4797 36552
rect 5224 36550 5342 36724
rect 4792 36486 5342 36550
rect 3013 36484 5342 36486
rect 3013 36476 4797 36484
rect 3013 36316 4797 36326
rect 5224 36316 5342 36484
rect 3013 36250 3018 36316
rect 4792 36250 5342 36316
rect 3013 36240 4797 36250
rect 3013 36080 4797 36090
rect 5224 36080 5342 36250
rect 3013 36014 3018 36080
rect 4792 36014 5342 36080
rect 3013 36004 4797 36014
rect 3013 35844 4797 35854
rect 3013 35778 3018 35844
rect 4792 35842 4797 35844
rect 5224 35842 5342 36014
rect 4792 35778 5342 35842
rect 3013 35776 5342 35778
rect 3013 35768 4797 35776
rect 3013 35608 4797 35618
rect 5224 35608 5342 35776
rect 3013 35542 3018 35608
rect 4792 35542 5342 35608
rect 3013 35532 4797 35542
rect 3013 35372 4797 35382
rect 5224 35372 5342 35542
rect 3013 35306 3018 35372
rect 4792 35306 5342 35372
rect 3013 35296 4797 35306
rect 3013 35136 4797 35146
rect 5224 35136 5342 35306
rect 3013 35070 3018 35136
rect 4792 35070 5342 35136
rect 3013 35060 4797 35070
rect 3013 34900 4797 34910
rect 5224 34900 5342 35070
rect 3013 34834 3018 34900
rect 4792 34834 5342 34900
rect 3013 34824 4797 34834
rect 3013 34664 4797 34674
rect 5224 34664 5342 34834
rect 3013 34598 3018 34664
rect 4792 34598 5342 34664
rect 3013 34588 4797 34598
rect 3013 34428 4797 34438
rect 5224 34428 5342 34598
rect 3013 34362 3018 34428
rect 4792 34362 5342 34428
rect 3013 34352 4797 34362
rect 3013 34192 4797 34202
rect 5224 34192 5342 34362
rect 3013 34126 3018 34192
rect 4792 34126 5342 34192
rect 3013 34116 4797 34126
rect 3013 33956 4797 33966
rect 5224 33956 5342 34126
rect 3013 33890 3018 33956
rect 4792 33890 5342 33956
rect 3013 33880 4797 33890
rect 3013 33720 4797 33730
rect 5224 33720 5342 33890
rect 3013 33654 3018 33720
rect 4792 33654 5342 33720
rect 3013 33644 4797 33654
rect 3013 33484 4797 33494
rect 3013 33418 3018 33484
rect 4792 33482 4797 33484
rect 5224 33482 5342 33654
rect 4792 33418 5342 33482
rect 3013 33416 5342 33418
rect 3013 33408 4797 33416
rect 3013 33248 4797 33258
rect 5224 33248 5342 33416
rect 3013 33182 3018 33248
rect 4792 33182 5342 33248
rect 3013 33172 4797 33182
rect 3013 33012 4797 33022
rect 5224 33012 5342 33182
rect 3013 32946 3018 33012
rect 4792 32946 5342 33012
rect 3013 32936 4797 32946
rect 3013 32776 4797 32786
rect 5224 32776 5342 32946
rect 3013 32710 3018 32776
rect 4792 32710 5342 32776
rect 3013 32700 4797 32710
rect 3013 32540 4797 32550
rect 3013 32474 3018 32540
rect 4792 32538 4797 32540
rect 5224 32538 5342 32710
rect 4792 32474 5342 32538
rect 3013 32472 5342 32474
rect 3013 32464 4797 32472
rect 3013 32304 4797 32314
rect 5224 32304 5342 32472
rect 3013 32238 3018 32304
rect 4792 32238 5342 32304
rect 3013 32228 4797 32238
rect 3013 32068 4797 32078
rect 5224 32068 5342 32238
rect 3013 32002 3018 32068
rect 4792 32002 5342 32068
rect 3013 31992 4797 32002
rect 3011 31832 4795 31842
rect 5224 31832 5342 32002
rect 3011 31766 3016 31832
rect 4790 31766 5342 31832
rect 3011 31756 4795 31766
rect 3013 31596 4797 31606
rect 5224 31596 5342 31766
rect 3013 31530 3018 31596
rect 4792 31530 5342 31596
rect 3013 31520 4797 31530
rect 3013 31360 4797 31370
rect 5224 31360 5342 31530
rect 3013 31294 3018 31360
rect 4792 31294 5342 31360
rect 3013 31284 4797 31294
rect 3013 31120 4797 31130
rect 5224 31120 5342 31294
rect 3013 31054 3018 31120
rect 4792 31060 5342 31120
rect 4792 31054 4797 31060
rect 3013 31050 4797 31054
rect 3018 31044 4792 31050
rect 5224 30950 5342 31060
rect 5332 29648 5342 30950
rect 5642 30950 5754 38168
rect 12392 38102 12992 43318
rect 23260 43240 23738 43860
rect 27086 43240 27492 43860
rect 23260 41038 27492 43240
rect 23242 40588 27492 41038
rect 12392 37306 12400 38102
rect 5642 29648 5652 30950
rect 12392 30490 12992 37306
rect 19672 40458 20138 40530
rect 20651 40460 23031 40470
rect 20651 40458 20656 40460
rect 19672 40440 20656 40458
rect 12382 29694 12392 30490
rect 12984 29694 12994 30490
rect 19672 29840 19796 40440
rect 19994 40398 20656 40440
rect 19994 40222 20138 40398
rect 20651 40396 20656 40398
rect 23026 40396 23031 40460
rect 20651 40386 23031 40396
rect 20651 40224 23031 40234
rect 20651 40222 20656 40224
rect 19994 40162 20656 40222
rect 19994 39988 20138 40162
rect 20651 40160 20656 40162
rect 23026 40160 23031 40224
rect 20651 40150 23031 40160
rect 20649 39988 23029 39998
rect 19994 39928 20654 39988
rect 19994 39750 20138 39928
rect 20649 39924 20654 39928
rect 23024 39924 23029 39988
rect 20649 39914 23029 39924
rect 20649 39752 23029 39762
rect 20649 39750 20654 39752
rect 19994 39690 20654 39750
rect 19994 39514 20138 39690
rect 20649 39688 20654 39690
rect 23024 39688 23029 39752
rect 20649 39678 23029 39688
rect 20651 39516 23031 39526
rect 20651 39514 20656 39516
rect 19994 39454 20656 39514
rect 19994 39274 20138 39454
rect 20651 39452 20656 39454
rect 23026 39452 23031 39516
rect 20651 39442 23031 39452
rect 20649 39278 23029 39288
rect 20649 39274 20654 39278
rect 19994 39214 20654 39274
rect 23024 39214 23029 39278
rect 19994 39038 20138 39214
rect 20649 39204 23029 39214
rect 20651 39042 23031 39052
rect 20651 39038 20656 39042
rect 19994 38978 20656 39038
rect 23026 38978 23031 39042
rect 19994 38806 20138 38978
rect 20651 38968 23031 38978
rect 20649 38810 23029 38820
rect 20649 38806 20654 38810
rect 19994 38746 20654 38806
rect 23024 38746 23029 38810
rect 19994 38570 20138 38746
rect 20649 38736 23029 38746
rect 20651 38570 23031 38580
rect 19994 38510 20656 38570
rect 19994 38332 20138 38510
rect 20651 38506 20656 38510
rect 23026 38506 23031 38570
rect 20651 38496 23031 38506
rect 20649 38334 23029 38344
rect 20649 38332 20654 38334
rect 19994 38272 20654 38332
rect 19994 38100 20138 38272
rect 20649 38270 20654 38272
rect 23024 38270 23029 38334
rect 20649 38260 23029 38270
rect 20649 38100 23029 38108
rect 19994 38098 23029 38100
rect 19994 38040 20654 38098
rect 19994 37862 20138 38040
rect 20649 38034 20654 38040
rect 23024 38034 23029 38098
rect 20649 38024 23029 38034
rect 20651 37862 23031 37872
rect 19994 37802 20656 37862
rect 19994 37624 20138 37802
rect 20651 37798 20656 37802
rect 23026 37798 23031 37862
rect 20651 37788 23031 37798
rect 20651 37626 23031 37636
rect 20651 37624 20656 37626
rect 19994 37564 20656 37624
rect 19994 37388 20138 37564
rect 20651 37562 20656 37564
rect 23026 37562 23031 37626
rect 20651 37552 23031 37562
rect 20651 37390 23031 37400
rect 20651 37388 20656 37390
rect 19994 37328 20656 37388
rect 19994 37156 20138 37328
rect 20651 37326 20656 37328
rect 23026 37326 23031 37390
rect 20651 37316 23031 37326
rect 20649 37156 23029 37166
rect 19994 37096 20654 37156
rect 19994 36918 20138 37096
rect 20649 37092 20654 37096
rect 23024 37092 23029 37156
rect 20649 37082 23029 37092
rect 20653 36920 23033 36930
rect 20653 36918 20658 36920
rect 19994 36858 20658 36918
rect 19994 36680 20138 36858
rect 20653 36856 20658 36858
rect 23028 36856 23033 36920
rect 20653 36846 23033 36856
rect 20651 36682 23031 36692
rect 20651 36680 20656 36682
rect 19994 36620 20656 36680
rect 19994 36442 20138 36620
rect 20651 36618 20656 36620
rect 23026 36618 23031 36682
rect 20651 36608 23031 36618
rect 20653 36446 23033 36456
rect 20653 36442 20658 36446
rect 19994 36382 20658 36442
rect 23028 36382 23033 36446
rect 19994 36208 20138 36382
rect 20653 36372 23033 36382
rect 20653 36210 23033 36220
rect 20653 36208 20658 36210
rect 19994 36148 20658 36208
rect 19994 35972 20138 36148
rect 20653 36146 20658 36148
rect 23028 36146 23033 36210
rect 20653 36136 23033 36146
rect 20653 35976 23033 35986
rect 20653 35972 20658 35976
rect 19994 35912 20658 35972
rect 23028 35912 23033 35976
rect 19994 35736 20138 35912
rect 20653 35902 23033 35912
rect 20649 35738 23029 35748
rect 20649 35736 20654 35738
rect 19994 35676 20654 35736
rect 19994 35498 20138 35676
rect 20649 35674 20654 35676
rect 23024 35674 23029 35738
rect 20649 35664 23029 35674
rect 20649 35500 23029 35510
rect 20649 35498 20654 35500
rect 19994 35438 20654 35498
rect 19994 35264 20138 35438
rect 20649 35436 20654 35438
rect 23024 35436 23029 35500
rect 20649 35426 23029 35436
rect 20651 35266 23031 35276
rect 20651 35264 20656 35266
rect 19994 35204 20656 35264
rect 19994 35030 20138 35204
rect 20651 35202 20656 35204
rect 23026 35202 23031 35266
rect 20651 35192 23031 35202
rect 20651 35030 23031 35040
rect 19994 34970 20656 35030
rect 19994 34792 20138 34970
rect 20651 34966 20656 34970
rect 23026 34966 23031 35030
rect 20651 34956 23031 34966
rect 20653 34794 23033 34804
rect 20653 34792 20658 34794
rect 19994 34732 20658 34792
rect 19994 34558 20138 34732
rect 20653 34730 20658 34732
rect 23028 34730 23033 34794
rect 20653 34720 23033 34730
rect 20649 34560 23029 34570
rect 20649 34558 20654 34560
rect 19994 34498 20654 34558
rect 19994 34320 20138 34498
rect 20649 34496 20654 34498
rect 23024 34496 23029 34560
rect 20649 34486 23029 34496
rect 20649 34322 23029 34332
rect 20649 34320 20654 34322
rect 19994 34260 20654 34320
rect 19994 34086 20138 34260
rect 20649 34258 20654 34260
rect 23024 34258 23029 34322
rect 20649 34248 23029 34258
rect 20651 34088 23031 34098
rect 20651 34086 20656 34088
rect 19994 34026 20656 34086
rect 19994 33846 20138 34026
rect 20651 34024 20656 34026
rect 23026 34024 23031 34088
rect 20651 34014 23031 34024
rect 20651 33850 23031 33860
rect 20651 33846 20656 33850
rect 19994 33786 20656 33846
rect 23026 33786 23031 33850
rect 19994 33614 20138 33786
rect 20651 33776 23031 33786
rect 20651 33614 23031 33624
rect 19994 33554 20656 33614
rect 19994 33380 20138 33554
rect 20651 33550 20656 33554
rect 23026 33550 23031 33614
rect 20651 33540 23031 33550
rect 20651 33380 23031 33390
rect 19994 33320 20656 33380
rect 19994 33142 20138 33320
rect 20651 33316 20656 33320
rect 23026 33316 23031 33380
rect 20651 33306 23031 33316
rect 20651 33144 23031 33154
rect 20651 33142 20656 33144
rect 19994 33082 20656 33142
rect 19994 32904 20138 33082
rect 20651 33080 20656 33082
rect 23026 33080 23031 33144
rect 20651 33070 23031 33080
rect 20651 32906 23031 32916
rect 20651 32904 20656 32906
rect 19994 32844 20656 32904
rect 19994 32670 20138 32844
rect 20651 32842 20656 32844
rect 23026 32842 23031 32906
rect 20651 32832 23031 32842
rect 20653 32672 23033 32682
rect 20653 32670 20658 32672
rect 19994 32610 20658 32670
rect 19994 32438 20138 32610
rect 20653 32608 20658 32610
rect 23028 32608 23033 32672
rect 20653 32598 23033 32608
rect 20653 32438 23033 32448
rect 19994 32378 20658 32438
rect 19994 32196 20138 32378
rect 20653 32374 20658 32378
rect 23028 32374 23033 32438
rect 20653 32364 23033 32374
rect 20651 32198 23031 32208
rect 20651 32196 20656 32198
rect 19994 32136 20656 32196
rect 19994 31962 20138 32136
rect 20651 32134 20656 32136
rect 23026 32134 23031 32198
rect 20651 32124 23031 32134
rect 20651 31964 23031 31974
rect 20651 31962 20656 31964
rect 19994 31902 20656 31962
rect 19994 31724 20138 31902
rect 20651 31900 20656 31902
rect 23026 31900 23031 31964
rect 20651 31890 23031 31900
rect 20651 31726 23031 31736
rect 20651 31724 20656 31726
rect 19994 31664 20656 31724
rect 19994 31490 20138 31664
rect 20651 31662 20656 31664
rect 23026 31662 23031 31726
rect 20651 31652 23031 31662
rect 20651 31492 23031 31502
rect 20651 31490 20656 31492
rect 19994 31430 20656 31490
rect 19994 31254 20138 31430
rect 20651 31428 20656 31430
rect 23026 31428 23031 31492
rect 20651 31418 23031 31428
rect 20651 31256 23031 31266
rect 20651 31254 20656 31256
rect 19994 31194 20656 31254
rect 19994 31018 20138 31194
rect 20651 31192 20656 31194
rect 23026 31192 23031 31256
rect 20651 31182 23031 31192
rect 20649 31020 23029 31030
rect 20649 31018 20654 31020
rect 19994 30958 20654 31018
rect 19994 30780 20138 30958
rect 20649 30956 20654 30958
rect 23024 30956 23029 31020
rect 20649 30946 23029 30956
rect 20651 30782 23031 30792
rect 20651 30780 20656 30782
rect 19994 30720 20656 30780
rect 19994 30544 20138 30720
rect 20651 30718 20656 30720
rect 23026 30718 23031 30782
rect 20651 30708 23031 30718
rect 20651 30546 23031 30556
rect 20651 30544 20656 30546
rect 19994 30484 20656 30544
rect 19994 30308 20138 30484
rect 20651 30482 20656 30484
rect 23026 30482 23031 30546
rect 20651 30472 23031 30482
rect 20651 30312 23031 30322
rect 20651 30308 20656 30312
rect 19994 30248 20656 30308
rect 23026 30248 23031 30312
rect 19994 30070 20138 30248
rect 20651 30238 23031 30248
rect 20651 30074 23031 30084
rect 20651 30070 20656 30074
rect 19994 30010 20656 30070
rect 23026 30010 23031 30074
rect 19994 29840 20138 30010
rect 20651 30000 23031 30010
rect 19672 29836 20138 29840
rect 20653 29840 23033 29850
rect 20653 29836 20658 29840
rect 19672 29776 20658 29836
rect 23028 29776 23033 29840
rect 12400 22914 12992 29694
rect 19672 29634 20138 29776
rect 20653 29766 23033 29776
rect 23242 27192 25116 40588
rect 21049 25056 23029 25066
rect 21049 24992 21054 25056
rect 23024 25054 23029 25056
rect 23241 25054 25116 27192
rect 23024 24994 25116 25054
rect 23024 24992 23029 24994
rect 21049 24982 23029 24992
rect 21049 24700 23029 24710
rect 21049 24636 21054 24700
rect 23024 24698 23029 24700
rect 23241 24698 25116 24994
rect 23024 24638 25116 24698
rect 23024 24636 23029 24638
rect 21049 24626 23029 24636
rect 21049 24342 23029 24352
rect 21049 24278 21054 24342
rect 23024 24340 23029 24342
rect 23241 24340 25116 24638
rect 23024 24280 25116 24340
rect 23024 24278 23029 24280
rect 21049 24268 23029 24278
rect 21049 23986 23029 23996
rect 21049 23922 21054 23986
rect 23024 23984 23029 23986
rect 23241 23984 25116 24280
rect 23024 23924 25116 23984
rect 23024 23922 23029 23924
rect 21049 23912 23029 23922
rect 21047 23632 23027 23642
rect 21047 23568 21052 23632
rect 23022 23630 23027 23632
rect 23241 23630 25116 23924
rect 23022 23570 25116 23630
rect 23022 23568 23027 23570
rect 21047 23558 23027 23568
rect 21049 23274 23029 23284
rect 21049 23210 21054 23274
rect 23024 23272 23029 23274
rect 23241 23272 25116 23570
rect 23024 23212 25116 23272
rect 23024 23210 23029 23212
rect 21049 23200 23029 23210
rect 21049 22920 23029 22930
rect 21049 22856 21054 22920
rect 23024 22918 23029 22920
rect 23241 22918 25116 23212
rect 23024 22858 25116 22918
rect 23024 22856 23029 22858
rect 21049 22846 23029 22856
rect 19804 22772 19984 22777
rect 18468 22684 18992 22689
rect 18468 22294 18478 22684
rect 18982 22294 18992 22684
rect 19804 22660 19814 22772
rect 19974 22660 19984 22772
rect 19804 22655 19984 22660
rect 21049 22562 23029 22572
rect 21049 22498 21054 22562
rect 23024 22560 23029 22562
rect 23241 22560 25116 22858
rect 23024 22500 25116 22560
rect 23024 22498 23029 22500
rect 21049 22488 23029 22498
rect 18468 22289 18992 22294
rect 21049 22206 23029 22216
rect 21049 22142 21054 22206
rect 23024 22204 23029 22206
rect 23241 22204 25116 22500
rect 23024 22144 25116 22204
rect 23024 22142 23029 22144
rect 21049 22132 23029 22142
rect 12400 22072 12992 22118
rect 4775 15710 6573 15720
rect 4775 15648 4780 15710
rect 6568 15708 6573 15710
rect 7246 15708 7796 22040
rect 21049 21852 23029 21862
rect 21049 21788 21054 21852
rect 23024 21850 23029 21852
rect 23241 21850 25116 22144
rect 23024 21790 25116 21850
rect 23024 21788 23029 21790
rect 21049 21778 23029 21788
rect 21049 21494 23029 21504
rect 21049 21430 21054 21494
rect 23024 21492 23029 21494
rect 23241 21492 25116 21790
rect 23024 21432 25116 21492
rect 23024 21430 23029 21432
rect 21049 21420 23029 21430
rect 19800 21144 19980 21149
rect 19800 21030 19810 21144
rect 19970 21030 19980 21144
rect 21049 21140 23029 21150
rect 21049 21076 21054 21140
rect 23024 21138 23029 21140
rect 23241 21138 25116 21432
rect 23024 21078 25116 21138
rect 23024 21076 23029 21078
rect 21049 21066 23029 21076
rect 19800 21025 19980 21030
rect 21047 20782 23027 20792
rect 21047 20718 21052 20782
rect 23022 20780 23027 20782
rect 23241 20780 25116 21078
rect 23022 20720 25116 20780
rect 23022 20718 23027 20720
rect 21047 20708 23027 20718
rect 6568 15648 7796 15708
rect 4775 15646 7796 15648
rect 4775 15638 6573 15646
rect 4775 15474 6573 15484
rect 4775 15412 4780 15474
rect 6568 15472 6794 15474
rect 7246 15472 7796 15646
rect 6568 15412 7796 15472
rect 4775 15410 7796 15412
rect 4775 15402 6573 15410
rect 4775 15238 6573 15248
rect 4775 15176 4780 15238
rect 6568 15236 6794 15238
rect 7246 15236 7796 15410
rect 6568 15176 7796 15236
rect 4775 15174 7796 15176
rect 4775 15166 6573 15174
rect 4775 15002 6573 15012
rect 7246 15002 7796 15174
rect 4775 14940 4780 15002
rect 6568 14940 7796 15002
rect 4775 14930 6573 14940
rect 4775 14768 6573 14776
rect 4775 14766 6794 14768
rect 7246 14766 7796 14940
rect 4775 14704 4780 14766
rect 6568 14704 7796 14766
rect 4775 14694 6573 14704
rect 4775 14530 6573 14540
rect 7246 14530 7796 14704
rect 4775 14468 4780 14530
rect 6568 14468 7796 14530
rect 4775 14458 6573 14468
rect 4775 14294 6573 14304
rect 7246 14294 7796 14468
rect 4775 14232 4780 14294
rect 6568 14232 7796 14294
rect 4775 14230 6794 14232
rect 4775 14222 6573 14230
rect 4775 14058 6573 14068
rect 7246 14058 7796 14232
rect 4775 13996 4780 14058
rect 6568 13996 7796 14058
rect 4775 13986 6573 13996
rect 4775 13824 6573 13832
rect 4775 13822 6794 13824
rect 7246 13822 7796 13996
rect 4775 13760 4780 13822
rect 6568 13760 7796 13822
rect 4775 13750 6573 13760
rect 4775 13586 6573 13596
rect 7246 13586 7796 13760
rect 4775 13524 4780 13586
rect 6568 13524 7796 13586
rect 4775 13514 6573 13524
rect 4775 13350 6573 13360
rect 7246 13350 7796 13524
rect 4775 13288 4780 13350
rect 6568 13288 7796 13350
rect 4775 13286 6794 13288
rect 4775 13278 6573 13286
rect 4775 13116 6573 13124
rect 7246 13116 7796 13288
rect 4775 13114 7796 13116
rect 4775 13052 4780 13114
rect 6568 13054 7796 13114
rect 6568 13052 6794 13054
rect 4775 13050 6794 13052
rect 4775 13042 6573 13050
rect 4775 12880 6573 12888
rect 7246 12880 7796 13054
rect 4775 12878 7796 12880
rect 4775 12816 4780 12878
rect 6568 12818 7796 12878
rect 6568 12816 6794 12818
rect 4775 12814 6794 12816
rect 4775 12806 6573 12814
rect 7246 12652 7796 12818
rect 9120 20558 19600 20600
rect 9120 20556 14540 20558
rect 9120 20486 9172 20556
rect 11540 20486 11808 20556
rect 14176 20488 14540 20556
rect 16908 20556 19600 20558
rect 16908 20488 17176 20556
rect 14176 20486 17176 20488
rect 19544 20486 19600 20556
rect 9120 20200 19600 20486
rect 21049 20424 23029 20434
rect 21049 20360 21054 20424
rect 23024 20422 23029 20424
rect 23241 20422 25116 20720
rect 23024 20362 25116 20422
rect 23024 20360 23029 20362
rect 21049 20350 23029 20360
rect 9120 20130 9172 20200
rect 11540 20130 11808 20200
rect 14176 20130 14540 20200
rect 16908 20130 17176 20200
rect 19544 20130 19600 20200
rect 9120 19844 19600 20130
rect 21047 20072 23027 20082
rect 21047 20008 21052 20072
rect 23022 20070 23027 20072
rect 23241 20070 25116 20362
rect 23022 20010 25116 20070
rect 23022 20008 23027 20010
rect 21047 19998 23027 20008
rect 9120 19774 9172 19844
rect 11540 19774 11808 19844
rect 14176 19774 14540 19844
rect 16908 19774 17176 19844
rect 19544 19774 19600 19844
rect 9120 19490 19600 19774
rect 21049 19714 23029 19724
rect 21049 19650 21054 19714
rect 23024 19712 23029 19714
rect 23241 19712 25116 20010
rect 23024 19652 25116 19712
rect 23024 19650 23029 19652
rect 21049 19640 23029 19650
rect 9120 19420 9172 19490
rect 11540 19488 19600 19490
rect 11540 19420 11808 19488
rect 9120 19418 11808 19420
rect 14176 19486 19600 19488
rect 14176 19418 14540 19486
rect 9120 19416 14540 19418
rect 16908 19416 17176 19486
rect 19544 19416 19600 19486
rect 9120 19132 19600 19416
rect 21047 19360 23027 19370
rect 21047 19296 21052 19360
rect 23022 19358 23027 19360
rect 23241 19358 25116 19652
rect 23022 19298 25116 19358
rect 23022 19296 23027 19298
rect 21047 19286 23027 19296
rect 9120 19062 9172 19132
rect 11540 19062 11808 19132
rect 14176 19062 14540 19132
rect 16908 19062 17176 19132
rect 19544 19062 19600 19132
rect 9120 18776 19600 19062
rect 21049 19002 23029 19012
rect 21049 18938 21054 19002
rect 23024 19000 23029 19002
rect 23241 19000 25116 19298
rect 23024 18940 25116 19000
rect 23024 18938 23029 18940
rect 21049 18928 23029 18938
rect 9120 18706 9172 18776
rect 11540 18706 11808 18776
rect 14176 18706 14540 18776
rect 16908 18706 17176 18776
rect 19544 18706 19600 18776
rect 9120 18420 19600 18706
rect 21047 18646 23027 18656
rect 21047 18582 21052 18646
rect 23022 18644 23027 18646
rect 23241 18644 25116 18940
rect 23022 18584 25116 18644
rect 23022 18582 23027 18584
rect 21047 18572 23027 18582
rect 9120 18350 9172 18420
rect 11540 18350 11808 18420
rect 14176 18350 14540 18420
rect 16908 18350 17176 18420
rect 19544 18350 19600 18420
rect 9120 18064 19600 18350
rect 21049 18290 23029 18300
rect 21049 18226 21054 18290
rect 23024 18288 23029 18290
rect 23241 18288 25116 18584
rect 23024 18228 25116 18288
rect 23024 18226 23029 18228
rect 21049 18216 23029 18226
rect 9120 17994 9172 18064
rect 11540 17994 11808 18064
rect 14176 17994 14540 18064
rect 16908 17994 17176 18064
rect 19544 17994 19600 18064
rect 9120 17708 19600 17994
rect 21049 17934 23029 17944
rect 21049 17870 21054 17934
rect 23024 17932 23029 17934
rect 23241 17932 25116 18228
rect 23024 17872 25116 17932
rect 23024 17870 23029 17872
rect 21049 17860 23029 17870
rect 9120 17638 9172 17708
rect 11540 17638 11808 17708
rect 14176 17638 14540 17708
rect 16908 17706 19600 17708
rect 16908 17638 17176 17706
rect 9120 17636 17176 17638
rect 19544 17636 19600 17706
rect 9120 17352 19600 17636
rect 21049 17578 23029 17588
rect 21049 17514 21054 17578
rect 23024 17576 23029 17578
rect 23241 17576 25116 17872
rect 23024 17516 25116 17576
rect 23024 17514 23029 17516
rect 21049 17504 23029 17514
rect 9120 17282 9172 17352
rect 11540 17282 11808 17352
rect 14176 17282 14540 17352
rect 16908 17282 17176 17352
rect 19544 17282 19600 17352
rect 9120 16996 19600 17282
rect 21049 17222 23029 17232
rect 21049 17158 21054 17222
rect 23024 17220 23029 17222
rect 23241 17220 25116 17516
rect 23024 17160 25116 17220
rect 23024 17158 23029 17160
rect 21049 17148 23029 17158
rect 9120 16926 9172 16996
rect 11540 16926 11808 16996
rect 14176 16926 14540 16996
rect 16908 16926 17176 16996
rect 19544 16926 19600 16996
rect 9120 16640 19600 16926
rect 21049 16866 23029 16876
rect 21049 16802 21054 16866
rect 23024 16864 23029 16866
rect 23241 16864 25116 17160
rect 23024 16804 25116 16864
rect 23024 16802 23029 16804
rect 21049 16792 23029 16802
rect 9120 16570 9172 16640
rect 11540 16570 11808 16640
rect 14176 16570 14540 16640
rect 16908 16570 17176 16640
rect 19544 16570 19600 16640
rect 9120 16286 19600 16570
rect 21047 16510 23027 16520
rect 21047 16446 21052 16510
rect 23022 16508 23027 16510
rect 23241 16508 25116 16804
rect 23022 16448 25116 16508
rect 23022 16446 23027 16448
rect 21047 16436 23027 16446
rect 9120 16284 11808 16286
rect 9120 16214 9172 16284
rect 11540 16216 11808 16284
rect 14176 16284 19600 16286
rect 14176 16216 14540 16284
rect 11540 16214 14540 16216
rect 16908 16214 17176 16284
rect 19544 16214 19600 16284
rect 9120 15928 19600 16214
rect 21049 16154 23029 16164
rect 21049 16090 21054 16154
rect 23024 16152 23029 16154
rect 23241 16152 25116 16448
rect 23024 16092 25116 16152
rect 23024 16090 23029 16092
rect 21049 16080 23029 16090
rect 9120 15858 9172 15928
rect 11540 15858 11808 15928
rect 14176 15926 17176 15928
rect 14176 15858 14540 15926
rect 9120 15856 14540 15858
rect 16908 15858 17176 15926
rect 19544 15858 19600 15928
rect 16908 15856 19600 15858
rect 9120 15572 19600 15856
rect 21049 15800 23029 15810
rect 21049 15736 21054 15800
rect 23024 15798 23029 15800
rect 23241 15798 25116 16092
rect 23024 15738 25116 15798
rect 23024 15736 23029 15738
rect 21049 15726 23029 15736
rect 9120 15502 9172 15572
rect 11540 15502 11808 15572
rect 14176 15502 14540 15572
rect 16908 15502 17176 15572
rect 19544 15502 19600 15572
rect 9120 15216 19600 15502
rect 21049 15442 23029 15452
rect 21049 15378 21054 15442
rect 23024 15440 23029 15442
rect 23241 15440 25116 15738
rect 23024 15380 25116 15440
rect 23024 15378 23029 15380
rect 21049 15368 23029 15378
rect 9120 15146 9172 15216
rect 11540 15146 11808 15216
rect 14176 15146 14540 15216
rect 16908 15146 17176 15216
rect 19544 15146 19600 15216
rect 9120 14860 19600 15146
rect 21049 15086 23029 15096
rect 21049 15022 21054 15086
rect 23024 15084 23029 15086
rect 23241 15084 25116 15380
rect 23024 15024 25116 15084
rect 23024 15022 23029 15024
rect 21049 15012 23029 15022
rect 9120 14790 9172 14860
rect 11540 14790 11808 14860
rect 14176 14790 14540 14860
rect 16908 14790 17176 14860
rect 19544 14790 19600 14860
rect 9120 14504 19600 14790
rect 21049 14732 23029 14742
rect 23241 14732 25116 15024
rect 21049 14668 21054 14732
rect 23024 14672 25116 14732
rect 23024 14668 23029 14672
rect 21049 14658 23029 14668
rect 9120 14434 9172 14504
rect 11540 14434 11808 14504
rect 14176 14434 14540 14504
rect 16908 14434 17176 14504
rect 19544 14434 19600 14504
rect 9120 14148 19600 14434
rect 21049 14374 23029 14384
rect 21049 14310 21054 14374
rect 23024 14372 23029 14374
rect 23241 14372 25116 14672
rect 23024 14312 25116 14372
rect 23024 14310 23029 14312
rect 21049 14300 23029 14310
rect 9120 14078 9172 14148
rect 11540 14078 11808 14148
rect 14176 14146 17176 14148
rect 14176 14078 14540 14146
rect 9120 14076 14540 14078
rect 16908 14078 17176 14146
rect 19544 14078 19600 14148
rect 16908 14076 19600 14078
rect 9120 13792 19600 14076
rect 9120 13722 9172 13792
rect 11540 13722 11808 13792
rect 14176 13722 14540 13792
rect 16908 13722 17176 13792
rect 19544 13722 19600 13792
rect 9120 13436 19600 13722
rect 21047 13790 23029 13798
rect 23241 13790 25116 14312
rect 21047 13788 25116 13790
rect 21047 13730 21052 13788
rect 23024 13730 25116 13788
rect 21047 13728 25116 13730
rect 21047 13720 23029 13728
rect 9120 13366 9172 13436
rect 11540 13366 11808 13436
rect 14176 13366 14540 13436
rect 16908 13366 17176 13436
rect 19544 13366 19600 13436
rect 9120 13080 19600 13366
rect 21047 13436 23029 13442
rect 23241 13436 25116 13728
rect 21047 13432 25116 13436
rect 21047 13374 21052 13432
rect 23024 13374 25116 13432
rect 21047 13364 23029 13374
rect 9120 13010 9172 13080
rect 11540 13010 11808 13080
rect 14176 13010 14540 13080
rect 16908 13010 17176 13080
rect 19544 13010 19600 13080
rect 9120 12724 19600 13010
rect 21047 13078 23029 13086
rect 23241 13078 25116 13374
rect 21047 13076 25116 13078
rect 21047 13018 21052 13076
rect 23024 13018 25116 13076
rect 21047 13016 25116 13018
rect 21047 13008 23029 13016
rect 9120 12654 9172 12724
rect 11540 12654 11808 12724
rect 14176 12654 14540 12724
rect 16908 12654 17176 12724
rect 19544 12654 19600 12724
rect 9120 12652 19600 12654
rect 21047 12722 23029 12730
rect 23241 12722 25116 13016
rect 21047 12720 25116 12722
rect 21047 12662 21052 12720
rect 23024 12662 25116 12720
rect 21047 12660 25116 12662
rect 21047 12652 23029 12660
rect 4768 12642 19600 12652
rect 4768 12580 4780 12642
rect 6568 12580 19600 12642
rect 4768 12406 19600 12580
rect 4768 12344 4780 12406
rect 6568 12368 19600 12406
rect 6568 12344 9172 12368
rect 4768 12298 9172 12344
rect 11540 12298 11808 12368
rect 14176 12298 14540 12368
rect 16908 12298 17178 12368
rect 19546 12298 19600 12368
rect 4768 12170 19600 12298
rect 21047 12366 23029 12374
rect 23241 12366 25116 12660
rect 21047 12364 25116 12366
rect 21047 12306 21052 12364
rect 23024 12306 25116 12364
rect 21047 12304 25116 12306
rect 21047 12296 23029 12304
rect 4768 12108 4780 12170
rect 6568 12108 19600 12170
rect 4768 12012 19600 12108
rect 4768 11942 9172 12012
rect 11540 11942 11808 12012
rect 14176 11942 14540 12012
rect 16908 11942 17178 12012
rect 19546 11942 19600 12012
rect 4768 11934 19600 11942
rect 21047 12010 23029 12018
rect 23241 12010 25116 12304
rect 21047 12008 25116 12010
rect 21047 11950 21052 12008
rect 23024 11950 25116 12008
rect 21047 11948 25116 11950
rect 21047 11940 23029 11948
rect 4768 11872 4780 11934
rect 6568 11872 19600 11934
rect 4768 11698 19600 11872
rect 4768 11636 4780 11698
rect 6568 11656 19600 11698
rect 6568 11646 9170 11656
rect 6568 11636 7796 11646
rect 4768 11628 7796 11636
rect 4775 11626 6573 11628
rect 4775 11464 6573 11472
rect 4775 11462 6794 11464
rect 4775 11400 4780 11462
rect 6568 11460 6794 11462
rect 7246 11460 7796 11628
rect 6568 11400 7796 11460
rect 4775 11398 7796 11400
rect 4775 11390 6573 11398
rect 4775 11226 6573 11236
rect 4775 11164 4780 11226
rect 6568 11224 6794 11226
rect 7246 11224 7796 11398
rect 6568 11164 7796 11224
rect 4775 11162 7796 11164
rect 4775 11154 6573 11162
rect 4775 10992 6573 11000
rect 4775 10990 6794 10992
rect 4775 10928 4780 10990
rect 6568 10988 6794 10990
rect 7246 10988 7796 11162
rect 6568 10928 7796 10988
rect 4775 10926 7796 10928
rect 4775 10918 6573 10926
rect 4775 10756 6573 10764
rect 4775 10754 6794 10756
rect 7246 10754 7796 10926
rect 4775 10692 4780 10754
rect 6568 10692 7796 10754
rect 4775 10682 6573 10692
rect 4775 10522 6573 10528
rect 4775 10518 6794 10522
rect 7246 10518 7796 10692
rect 4775 10456 4780 10518
rect 6568 10456 7796 10518
rect 4775 10446 6573 10456
rect 4775 10284 6573 10292
rect 4775 10282 6794 10284
rect 4775 10220 4780 10282
rect 6568 10280 6794 10282
rect 7246 10280 7796 10456
rect 6568 10220 7796 10280
rect 4775 10218 7796 10220
rect 4775 10210 6573 10218
rect 4775 10048 6573 10056
rect 4775 10046 6794 10048
rect 7246 10046 7796 10218
rect 4775 9984 4780 10046
rect 6568 9984 7796 10046
rect 4775 9974 6573 9984
rect 4775 9812 6573 9820
rect 4775 9810 6794 9812
rect 7246 9810 7796 9984
rect 4775 9748 4780 9810
rect 6568 9748 7796 9810
rect 4775 9738 6573 9748
rect 4775 9576 6573 9584
rect 4775 9574 6794 9576
rect 7246 9574 7796 9748
rect 4775 9512 4780 9574
rect 6568 9512 7796 9574
rect 4775 9502 6573 9512
rect 4775 9338 6573 9348
rect 7246 9338 7796 9512
rect 4775 9276 4780 9338
rect 6568 9276 7796 9338
rect 4775 9274 6794 9276
rect 4775 9266 6573 9274
rect 4775 9102 6573 9112
rect 4775 9038 4780 9102
rect 6568 9100 6573 9102
rect 6568 9098 6794 9100
rect 7246 9098 7796 9276
rect 6568 9038 7796 9098
rect 4775 9036 7796 9038
rect 4775 9028 6573 9036
rect 4775 8868 6573 8878
rect 7246 8868 7796 9036
rect 4775 8804 4780 8868
rect 6568 8806 7796 8868
rect 6568 8804 6794 8806
rect 4775 8794 6573 8804
rect 4775 8632 6573 8642
rect 4775 8568 4780 8632
rect 6568 8630 6794 8632
rect 7246 8630 7796 8806
rect 6568 8568 7796 8630
rect 4775 8558 6573 8568
rect 7246 2800 7796 8568
rect 9120 11586 9170 11646
rect 11538 11586 11808 11656
rect 14176 11586 14540 11656
rect 16908 11586 17176 11656
rect 19544 11586 19600 11656
rect 9120 11300 19600 11586
rect 21047 11656 23029 11662
rect 23241 11656 25116 11948
rect 21047 11652 25116 11656
rect 21047 11594 21052 11652
rect 23024 11594 25116 11652
rect 21047 11584 23029 11594
rect 9120 11230 9170 11300
rect 11538 11230 11808 11300
rect 14176 11230 14540 11300
rect 16908 11230 17176 11300
rect 19544 11230 19600 11300
rect 9120 10946 19600 11230
rect 21047 11300 23029 11306
rect 23241 11300 25116 11594
rect 21047 11296 25116 11300
rect 21047 11238 21052 11296
rect 23024 11238 25116 11296
rect 21047 11228 23029 11238
rect 9120 10944 14540 10946
rect 9120 10874 9170 10944
rect 11538 10874 11808 10944
rect 14176 10876 14540 10944
rect 16908 10944 19600 10946
rect 16908 10876 17176 10944
rect 14176 10874 17176 10876
rect 19544 10874 19600 10944
rect 9120 10588 19600 10874
rect 21047 10942 23029 10950
rect 23241 10942 25116 11238
rect 21047 10940 25116 10942
rect 21047 10882 21052 10940
rect 23024 10882 25116 10940
rect 21047 10880 25116 10882
rect 21047 10872 23029 10880
rect 9120 10518 9170 10588
rect 11538 10518 11808 10588
rect 14176 10586 17176 10588
rect 14176 10518 14538 10586
rect 9120 10516 14538 10518
rect 16906 10518 17176 10586
rect 19544 10518 19600 10588
rect 16906 10516 19600 10518
rect 21047 10586 23029 10594
rect 23241 10586 25116 10880
rect 21047 10584 25116 10586
rect 21047 10526 21052 10584
rect 23024 10526 25116 10584
rect 21047 10524 25116 10526
rect 21047 10516 23029 10524
rect 9120 10232 19600 10516
rect 9120 10162 9170 10232
rect 11538 10162 11808 10232
rect 14176 10162 14540 10232
rect 16908 10162 17176 10232
rect 19544 10162 19600 10232
rect 9120 9876 19600 10162
rect 21047 10230 23029 10238
rect 23241 10230 25116 10524
rect 21047 10228 25116 10230
rect 21047 10170 21052 10228
rect 23024 10170 25116 10228
rect 21047 10168 25116 10170
rect 21047 10160 23029 10168
rect 9120 9806 9170 9876
rect 11538 9806 11808 9876
rect 14176 9806 14540 9876
rect 16908 9806 17176 9876
rect 19544 9806 19600 9876
rect 9120 9520 19600 9806
rect 21047 9876 23029 9882
rect 23241 9876 25116 10168
rect 21047 9872 25116 9876
rect 21047 9814 21052 9872
rect 23024 9814 25116 9872
rect 21047 9812 25116 9814
rect 21047 9804 23029 9812
rect 9120 9450 9172 9520
rect 11540 9450 11808 9520
rect 14176 9450 14538 9520
rect 16906 9450 17176 9520
rect 19544 9450 19600 9520
rect 9120 9164 19600 9450
rect 21047 9520 23029 9526
rect 23241 9520 25116 9812
rect 21047 9516 25116 9520
rect 21047 9458 21052 9516
rect 23024 9458 25116 9516
rect 21047 9456 25116 9458
rect 21047 9448 23029 9456
rect 9120 9094 9172 9164
rect 11540 9094 11810 9164
rect 14178 9094 14538 9164
rect 16906 9094 17176 9164
rect 19544 9094 19600 9164
rect 9120 8808 19600 9094
rect 21047 9164 23029 9170
rect 23241 9164 25116 9456
rect 21047 9160 25116 9164
rect 21047 9102 21052 9160
rect 23024 9102 25116 9160
rect 21047 9100 25116 9102
rect 21047 9092 23029 9100
rect 9120 8806 11810 8808
rect 9120 8736 9172 8806
rect 11540 8738 11810 8806
rect 14178 8806 17176 8808
rect 14178 8738 14538 8806
rect 11540 8736 14538 8738
rect 16906 8738 17176 8806
rect 19544 8738 19600 8808
rect 16906 8736 19600 8738
rect 21047 8808 23029 8814
rect 23241 8808 25116 9100
rect 21047 8804 25116 8808
rect 21047 8746 21052 8804
rect 23024 8746 25116 8804
rect 21047 8744 25116 8746
rect 21047 8736 23029 8744
rect 9120 8452 19600 8736
rect 9120 8382 9172 8452
rect 11540 8382 11808 8452
rect 14176 8382 14538 8452
rect 16906 8382 17176 8452
rect 19544 8382 19600 8452
rect 9120 8096 19600 8382
rect 21049 8452 23031 8458
rect 23241 8452 25116 8744
rect 21049 8448 25116 8452
rect 21049 8390 21054 8448
rect 23026 8390 25116 8448
rect 21049 8388 25116 8390
rect 21049 8380 23031 8388
rect 9120 8026 9172 8096
rect 11540 8026 11810 8096
rect 14178 8026 14540 8096
rect 16908 8026 17176 8096
rect 19544 8026 19600 8096
rect 9120 7742 19600 8026
rect 21047 8096 23029 8102
rect 23241 8096 25116 8388
rect 21047 8092 25116 8096
rect 21047 8034 21052 8092
rect 23024 8034 25116 8092
rect 21047 8032 25116 8034
rect 21047 8024 23029 8032
rect 9120 7740 14540 7742
rect 9120 7670 9172 7740
rect 11540 7670 11808 7740
rect 14176 7672 14540 7740
rect 16908 7740 19600 7742
rect 16908 7672 17176 7740
rect 14176 7670 17176 7672
rect 19544 7670 19600 7740
rect 9120 7384 19600 7670
rect 21047 7740 23029 7746
rect 23241 7740 25116 8032
rect 21047 7736 25116 7740
rect 21047 7678 21052 7736
rect 23024 7678 25116 7736
rect 21047 7676 25116 7678
rect 21047 7668 23029 7676
rect 9120 7314 9172 7384
rect 11540 7314 11808 7384
rect 14176 7314 14540 7384
rect 16908 7314 17176 7384
rect 19544 7314 19600 7384
rect 9120 7028 19600 7314
rect 21047 7384 23029 7390
rect 23241 7384 25116 7676
rect 21047 7380 25116 7384
rect 21047 7322 21052 7380
rect 23024 7322 25116 7380
rect 21047 7320 25116 7322
rect 21047 7312 23029 7320
rect 9120 6958 9172 7028
rect 11540 6958 11810 7028
rect 14178 7026 17176 7028
rect 14178 6958 14540 7026
rect 9120 6956 14540 6958
rect 16908 6958 17176 7026
rect 19544 6958 19600 7028
rect 16908 6956 19600 6958
rect 21047 7028 23029 7034
rect 23241 7028 25116 7320
rect 21047 7024 25116 7028
rect 21047 6966 21052 7024
rect 23024 6966 25116 7024
rect 21047 6964 25116 6966
rect 21047 6956 23029 6964
rect 9120 6672 19600 6956
rect 9120 6602 9172 6672
rect 11540 6602 11808 6672
rect 14176 6602 14540 6672
rect 16908 6602 17176 6672
rect 19544 6602 19600 6672
rect 9120 6316 19600 6602
rect 21047 6672 23029 6678
rect 23241 6672 25116 6964
rect 21047 6668 25116 6672
rect 21047 6610 21052 6668
rect 23024 6610 25116 6668
rect 21047 6608 25116 6610
rect 21047 6600 23029 6608
rect 9120 6246 9172 6316
rect 11540 6246 11810 6316
rect 14178 6246 14540 6316
rect 16908 6246 17176 6316
rect 19544 6246 19600 6316
rect 9120 5962 19600 6246
rect 21047 6316 23029 6322
rect 23241 6316 25116 6608
rect 21047 6312 25116 6316
rect 21047 6254 21052 6312
rect 23024 6254 25116 6312
rect 21047 6252 25116 6254
rect 21047 6244 23029 6252
rect 9120 5960 14540 5962
rect 9120 5890 9170 5960
rect 11538 5890 11810 5960
rect 14178 5892 14540 5960
rect 16908 5960 19600 5962
rect 16908 5892 17176 5960
rect 14178 5890 17176 5892
rect 19544 5890 19600 5960
rect 9120 5604 19600 5890
rect 21047 5960 23029 5966
rect 23241 5960 25116 6252
rect 21047 5956 25116 5960
rect 21047 5898 21052 5956
rect 23024 5898 25116 5956
rect 21047 5896 25116 5898
rect 21047 5888 23029 5896
rect 9120 5534 9172 5604
rect 11540 5534 11808 5604
rect 14176 5534 14540 5604
rect 16908 5534 17176 5604
rect 19544 5534 19600 5604
rect 9120 5248 19600 5534
rect 21047 5604 23029 5610
rect 23241 5604 25116 5896
rect 21047 5600 25116 5604
rect 21047 5542 21052 5600
rect 23024 5542 25116 5600
rect 21047 5540 25116 5542
rect 21047 5532 23029 5540
rect 9120 5246 11808 5248
rect 9120 5176 9172 5246
rect 11540 5178 11808 5246
rect 14176 5246 17176 5248
rect 14176 5178 14540 5246
rect 11540 5176 14540 5178
rect 16908 5178 17176 5246
rect 19544 5178 19600 5248
rect 16908 5176 19600 5178
rect 21047 5248 23029 5254
rect 23241 5248 25116 5540
rect 21047 5244 25116 5248
rect 21047 5186 21052 5244
rect 23024 5186 25116 5244
rect 21047 5184 25116 5186
rect 21047 5176 23029 5184
rect 9120 4892 19600 5176
rect 9120 4822 9172 4892
rect 11540 4822 11808 4892
rect 14176 4822 14540 4892
rect 16908 4822 17176 4892
rect 19544 4822 19600 4892
rect 9120 4536 19600 4822
rect 21047 4892 23029 4898
rect 23241 4892 25116 5184
rect 21047 4888 25116 4892
rect 21047 4830 21052 4888
rect 23024 4830 25116 4888
rect 21047 4828 25116 4830
rect 21047 4820 23029 4828
rect 9120 4466 9172 4536
rect 11540 4466 11808 4536
rect 14176 4466 14540 4536
rect 16908 4466 17176 4536
rect 19544 4466 19600 4536
rect 9120 4180 19600 4466
rect 21047 4536 23029 4542
rect 23241 4536 25116 4828
rect 21047 4532 25116 4536
rect 21047 4474 21052 4532
rect 23024 4474 25116 4532
rect 21047 4472 25116 4474
rect 21047 4464 23029 4472
rect 9120 4110 9172 4180
rect 11540 4110 11808 4180
rect 14176 4110 14540 4180
rect 16908 4110 17176 4180
rect 19544 4110 19600 4180
rect 9120 3824 19600 4110
rect 21047 4180 23029 4186
rect 23241 4180 25116 4472
rect 21047 4176 25116 4180
rect 21047 4118 21052 4176
rect 23024 4118 25116 4176
rect 21047 4116 25116 4118
rect 21047 4108 23029 4116
rect 9120 3754 9172 3824
rect 11540 3754 11808 3824
rect 14176 3754 14540 3824
rect 16908 3754 17176 3824
rect 19544 3754 19600 3824
rect 9120 3468 19600 3754
rect 21047 3824 23029 3830
rect 23241 3824 25116 4116
rect 21047 3820 25116 3824
rect 21047 3762 21052 3820
rect 23024 3762 25116 3820
rect 21047 3760 25116 3762
rect 21047 3752 23029 3760
rect 9120 3398 9172 3468
rect 11540 3398 11808 3468
rect 14176 3466 17176 3468
rect 14176 3398 14540 3466
rect 9120 3396 14540 3398
rect 16908 3398 17176 3466
rect 19544 3398 19600 3468
rect 16908 3396 19600 3398
rect 21047 3468 23029 3474
rect 23241 3468 25116 3760
rect 21047 3464 25116 3468
rect 21047 3406 21052 3464
rect 23024 3406 25116 3464
rect 21047 3404 25116 3406
rect 21047 3396 23029 3404
rect 9120 3112 19600 3396
rect 23241 3290 25116 3404
rect 23006 3226 25116 3290
rect 9120 3042 9172 3112
rect 11540 3042 11808 3112
rect 14176 3042 14540 3112
rect 16908 3042 17176 3112
rect 19544 3042 19600 3112
rect 9120 3000 19600 3042
rect 21047 3112 23029 3118
rect 23241 3112 25116 3226
rect 21047 3108 25116 3112
rect 21047 3050 21052 3108
rect 23024 3050 25116 3108
rect 21047 3048 25116 3050
rect 21047 3040 23029 3048
rect 23241 2734 25116 3048
rect 25640 2734 27498 40588
rect 210 2496 590 2501
rect 210 1048 220 2496
rect 580 1048 590 2496
rect 11172 2286 12202 2291
rect 6232 2272 7262 2277
rect 6232 1280 6242 2272
rect 7252 1280 7262 2272
rect 11172 1294 11182 2286
rect 12192 1294 12202 2286
rect 11172 1289 12202 1294
rect 16514 2286 17544 2291
rect 16514 1294 16524 2286
rect 17534 1294 17544 2286
rect 23241 1960 27498 2734
rect 16514 1289 17544 1294
rect 6232 1275 7262 1280
rect 210 1043 590 1048
rect 23242 1000 27498 1960
rect 23260 998 27498 1000
<< via3 >>
rect 3018 38138 4792 38204
rect 3018 37902 4792 37968
rect 3018 37666 4792 37732
rect 3018 37430 4792 37496
rect 3018 37194 4792 37260
rect 3018 36958 4792 37024
rect 3018 36722 4792 36788
rect 3018 36486 4792 36552
rect 3018 36250 4792 36316
rect 3018 36014 4792 36080
rect 3018 35778 4792 35844
rect 3018 35542 4792 35608
rect 3018 35306 4792 35372
rect 3018 35070 4792 35136
rect 3018 34834 4792 34900
rect 3018 34598 4792 34664
rect 3018 34362 4792 34428
rect 3018 34126 4792 34192
rect 3018 33890 4792 33956
rect 3018 33654 4792 33720
rect 3018 33418 4792 33484
rect 3018 33182 4792 33248
rect 3018 32946 4792 33012
rect 3018 32710 4792 32776
rect 3018 32474 4792 32540
rect 3018 32238 4792 32304
rect 3018 32002 4792 32068
rect 3016 31766 4790 31832
rect 3018 31530 4792 31596
rect 3018 31294 4792 31360
rect 3018 31060 4792 31120
rect 3018 31054 4792 31060
rect 5342 29648 5642 38168
rect 23738 43240 27086 43860
rect 12400 37306 12992 38102
rect 12392 29694 12984 30490
rect 19796 29840 19994 40440
rect 12400 22118 12992 22914
rect 18478 22294 18982 22684
rect 19814 22660 19974 22772
rect 19810 21030 19970 21144
rect 220 1048 580 2496
rect 6242 1280 7252 2272
rect 11182 1294 12192 2286
rect 16524 1294 17534 2286
<< metal4 >>
rect 802 45036 29378 45152
rect 800 44812 29378 45036
rect 800 44152 1198 44812
rect 200 2496 600 44152
rect 200 1048 220 2496
rect 580 1048 600 2496
rect 200 1000 600 1048
rect 800 1000 1200 44152
rect 5196 43656 5800 44450
rect 19592 43656 20196 44450
rect 5196 42640 20196 43656
rect 23594 43860 27180 44812
rect 23594 43240 23738 43860
rect 27086 43240 27180 43860
rect 23594 43176 27178 43240
rect 3017 38204 4793 38205
rect 3017 38138 3018 38204
rect 4792 38144 5024 38204
rect 5196 38168 5800 42640
rect 19592 40440 20196 42640
rect 4792 38138 4793 38144
rect 3017 38137 4793 38138
rect 3017 37968 4793 37969
rect 3017 37902 3018 37968
rect 4792 37964 4793 37968
rect 4792 37904 5024 37964
rect 4792 37902 4793 37904
rect 3017 37901 4793 37902
rect 3017 37732 4793 37733
rect 3017 37666 3018 37732
rect 4792 37730 4793 37732
rect 4792 37670 5024 37730
rect 4792 37666 4793 37670
rect 3017 37665 4793 37666
rect 3017 37496 4793 37497
rect 3017 37430 3018 37496
rect 4792 37494 4793 37496
rect 4792 37434 5024 37494
rect 4792 37430 4793 37434
rect 3017 37429 4793 37430
rect 3017 37260 4793 37261
rect 3017 37194 3018 37260
rect 4792 37258 4793 37260
rect 4792 37198 5024 37258
rect 4792 37194 4793 37198
rect 3017 37193 4793 37194
rect 3017 37024 4793 37025
rect 3017 36958 3018 37024
rect 4792 37022 4793 37024
rect 4792 36962 5024 37022
rect 4792 36958 4793 36962
rect 3017 36957 4793 36958
rect 3017 36788 4793 36789
rect 3017 36722 3018 36788
rect 4792 36722 4793 36788
rect 3017 36721 4793 36722
rect 3017 36552 4793 36553
rect 3017 36486 3018 36552
rect 4792 36550 4793 36552
rect 4792 36490 5024 36550
rect 4792 36486 4793 36490
rect 3017 36485 4793 36486
rect 3017 36316 4793 36317
rect 3017 36250 3018 36316
rect 4792 36314 4793 36316
rect 4792 36254 5024 36314
rect 4792 36250 4793 36254
rect 3017 36249 4793 36250
rect 3017 36080 4793 36081
rect 3017 36014 3018 36080
rect 4792 36078 4793 36080
rect 4792 36018 5024 36078
rect 4792 36014 4793 36018
rect 3017 36013 4793 36014
rect 3017 35844 4793 35845
rect 3017 35778 3018 35844
rect 4792 35842 4793 35844
rect 4792 35782 5024 35842
rect 4792 35778 4793 35782
rect 3017 35777 4793 35778
rect 3017 35608 4793 35609
rect 3017 35542 3018 35608
rect 4792 35606 4793 35608
rect 4792 35546 5024 35606
rect 4792 35542 4793 35546
rect 3017 35541 4793 35542
rect 3017 35372 4793 35373
rect 3017 35306 3018 35372
rect 4792 35370 4793 35372
rect 4792 35310 5024 35370
rect 4792 35306 4793 35310
rect 3017 35305 4793 35306
rect 3017 35136 4793 35137
rect 3017 35070 3018 35136
rect 4792 35134 4793 35136
rect 4792 35074 5024 35134
rect 4792 35070 4793 35074
rect 3017 35069 4793 35070
rect 3017 34900 4793 34901
rect 3017 34834 3018 34900
rect 4792 34896 4793 34900
rect 4792 34836 5024 34896
rect 4792 34834 4793 34836
rect 3017 34833 4793 34834
rect 3017 34664 4793 34665
rect 3017 34598 3018 34664
rect 4792 34660 4793 34664
rect 4792 34600 5024 34660
rect 4792 34598 4793 34600
rect 3017 34597 4793 34598
rect 3017 34428 4793 34429
rect 3017 34362 3018 34428
rect 4792 34426 4793 34428
rect 4792 34366 5024 34426
rect 4792 34362 4793 34366
rect 3017 34361 4793 34362
rect 3017 34192 4793 34193
rect 3017 34126 3018 34192
rect 4792 34190 4793 34192
rect 4792 34130 5024 34190
rect 4792 34126 4793 34130
rect 3017 34125 4793 34126
rect 3017 33956 4793 33957
rect 3017 33890 3018 33956
rect 4792 33952 4793 33956
rect 4792 33892 5024 33952
rect 4792 33890 4793 33892
rect 3017 33889 4793 33890
rect 3017 33720 4793 33721
rect 3017 33654 3018 33720
rect 4792 33716 4793 33720
rect 4792 33656 5024 33716
rect 4792 33654 4793 33656
rect 3017 33653 4793 33654
rect 3017 33484 4793 33485
rect 3017 33418 3018 33484
rect 4792 33424 5024 33484
rect 4792 33418 4793 33424
rect 3017 33417 4793 33418
rect 3017 33248 4793 33249
rect 3017 33182 3018 33248
rect 4792 33246 4793 33248
rect 4792 33186 5024 33246
rect 4792 33182 4793 33186
rect 3017 33181 4793 33182
rect 3017 33012 4793 33013
rect 3017 32946 3018 33012
rect 4792 33010 4793 33012
rect 4792 32950 5024 33010
rect 4792 32946 4793 32950
rect 3017 32945 4793 32946
rect 3017 32776 4793 32777
rect 3017 32710 3018 32776
rect 4792 32774 4793 32776
rect 4792 32714 5024 32774
rect 4792 32710 4793 32714
rect 3017 32709 4793 32710
rect 3017 32540 4793 32541
rect 3017 32474 3018 32540
rect 4792 32538 4793 32540
rect 4792 32478 5024 32538
rect 4792 32474 4793 32478
rect 3017 32473 4793 32474
rect 3017 32304 4793 32305
rect 3017 32238 3018 32304
rect 4792 32302 4793 32304
rect 4792 32242 5024 32302
rect 4792 32238 4793 32242
rect 3017 32237 4793 32238
rect 3017 32068 4793 32069
rect 3017 32002 3018 32068
rect 4792 32066 4793 32068
rect 4792 32006 5024 32066
rect 4792 32002 4793 32006
rect 3017 32001 4793 32002
rect 3015 31832 4791 31833
rect 3015 31766 3016 31832
rect 4790 31830 4791 31832
rect 4790 31770 5024 31830
rect 4790 31766 4791 31770
rect 3015 31765 4791 31766
rect 3017 31596 4793 31597
rect 3017 31530 3018 31596
rect 4792 31594 4793 31596
rect 4792 31534 5024 31594
rect 4792 31530 4793 31534
rect 3017 31529 4793 31530
rect 3017 31360 4793 31361
rect 3017 31294 3018 31360
rect 4792 31358 4793 31360
rect 4792 31298 5024 31358
rect 4792 31294 4793 31298
rect 3017 31293 4793 31294
rect 3018 31121 5024 31122
rect 3017 31120 5024 31121
rect 3017 31054 3018 31120
rect 4792 31060 5024 31120
rect 4792 31054 4793 31060
rect 3017 31053 4793 31054
rect 5196 29648 5342 38168
rect 5642 34338 5800 38168
rect 6054 38102 19352 38168
rect 6054 37306 12400 38102
rect 12992 37306 19352 38102
rect 6054 37250 19352 37306
rect 5642 33322 19350 34338
rect 5642 29648 5800 33322
rect 12986 30566 19352 30568
rect 6054 30490 19352 30566
rect 6054 29694 12392 30490
rect 12984 29694 19352 30490
rect 6054 29650 19352 29694
rect 19592 29840 19796 40440
rect 19994 29840 20196 40440
rect 6054 29648 15722 29650
rect 5196 26668 5800 29648
rect 19592 28066 20196 29840
rect 19592 27068 29358 28066
rect 19592 26668 20196 27068
rect 5188 25652 20196 26668
rect 5196 23220 5800 25652
rect 19592 23254 20196 25652
rect 6054 22914 19348 22968
rect 6054 22118 12400 22914
rect 12992 22684 19348 22914
rect 12992 22294 18478 22684
rect 18982 22294 19348 22684
rect 12992 22118 19348 22294
rect 6054 22050 19348 22118
rect 19788 22772 19994 22784
rect 19788 22660 19814 22772
rect 19974 22660 19994 22772
rect 19788 21144 19994 22660
rect 19788 21030 19810 21144
rect 19970 21030 19994 21144
rect 19788 21020 19994 21030
rect 11181 2286 12193 2287
rect 6241 2272 7253 2273
rect 6241 1280 6242 2272
rect 7252 1280 7253 2272
rect 11181 1294 11182 2286
rect 12192 1294 12193 2286
rect 11181 1293 12193 1294
rect 16523 2286 17535 2287
rect 16523 1294 16524 2286
rect 17534 1954 17535 2286
rect 17534 1664 26690 1954
rect 17534 1294 17535 1664
rect 16523 1293 17535 1294
rect 6241 1279 7253 1280
rect 6642 670 6824 1279
rect 11584 1134 11766 1293
rect 11584 1128 20612 1134
rect 11584 838 22816 1128
rect 18770 670 18952 672
rect 6642 380 18952 670
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18952 380
rect 22634 0 22816 838
rect 26498 0 26678 1664
rect 28218 198 29354 27068
rect 30362 198 30542 200
rect 28218 0 30542 198
<< rmetal4 >>
rect 4793 36726 5024 36786
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_0
timestamp 1723380300
transform 0 -1 16300 -1 0 26036
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_1
timestamp 1723380300
transform 0 -1 9090 -1 0 26036
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_2
timestamp 1723380300
transform 0 -1 16286 -1 0 33636
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_3
timestamp 1723380300
transform 0 -1 16270 -1 0 41236
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_4
timestamp 1723380300
transform 0 -1 9102 -1 0 33636
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_5
timestamp 1723380300
transform 0 -1 9084 -1 0 41234
box -3186 -3040 3186 3040
use sky130_fd_pr__nfet_01v8_72JNYZ  sky130_fd_pr__nfet_01v8_72JNYZ_0
timestamp 1723380300
transform 0 -1 18682 1 0 21641
box -211 -1110 211 1110
use sky130_fd_pr__nfet_01v8_83M5YB  sky130_fd_pr__nfet_01v8_83M5YB_1
timestamp 1723380300
transform 0 -1 21842 1 0 35117
box -5477 -1410 5477 1410
use sky130_fd_pr__nfet_01v8_T4HZYF  sky130_fd_pr__nfet_01v8_T4HZYF_0
timestamp 1723380300
transform 0 -1 22038 1 0 8419
box -5685 -1210 5685 1210
use sky130_fd_pr__nfet_01v8_T4HZYF  sky130_fd_pr__nfet_01v8_T4HZYF_1
timestamp 1723380300
transform 0 -1 22038 1 0 19683
box -5685 -1210 5685 1210
use sky130_fd_pr__pfet_01v8_2EV7WZ  sky130_fd_pr__pfet_01v8_2EV7WZ_0
timestamp 1723380300
transform 0 -1 5675 1 0 8017
box -521 -1119 521 1119
use sky130_fd_pr__pfet_01v8_3WZJZZ  sky130_fd_pr__pfet_01v8_3WZJZZ_0
timestamp 1723380300
transform 0 -1 5675 1 0 12139
box -3707 -1119 3707 1119
use sky130_fd_pr__pfet_01v8_3WZJZZ  sky130_fd_pr__pfet_01v8_3WZJZZ_1
timestamp 1723380300
transform 0 -1 3905 1 0 34631
box -3707 -1119 3707 1119
use sky130_fd_pr__pfet_01v8_S7TZH4  sky130_fd_pr__pfet_01v8_S7TZH4_0
timestamp 1723380300
transform 0 -1 17041 1 0 11799
box -9067 -2737 9067 2737
use sky130_fd_pr__pfet_01v8_S7TZH4  sky130_fd_pr__pfet_01v8_S7TZH4_1
timestamp 1723380300
transform 0 -1 11673 1 0 11799
box -9067 -2737 9067 2737
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
rlabel metal2 2798 1298 3794 2302 7 vdd
rlabel via1 11182 1294 12192 2286 7 vin_n
rlabel via1 16524 1294 17534 2286 7 vin_p
rlabel metal3 23978 1282 24988 2274 7 vss
rlabel via1 6242 1280 7252 2272 7 iref
rlabel metal4 12174 42648 13184 43640 7 vout
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal tristate
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal tristate
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal tristate
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal tristate
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal tristate
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal tristate
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal tristate
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal tristate
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal tristate
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal tristate
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal tristate
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal tristate
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal tristate
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal tristate
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal tristate
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal tristate
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal tristate
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal tristate
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal tristate
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal tristate
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal tristate
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal tristate
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal tristate
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal tristate
flabel metal4 200 1000 600 44152 1 FreeSans 2 0 0 0 VDPWR
port 53 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 2 0 0 0 VGND
port 54 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
