magic
tech sky130A
magscale 1 2
timestamp 1723380300
<< error_p >>
rect -324 981 -266 987
rect -206 981 -148 987
rect -88 981 -30 987
rect 30 981 88 987
rect 148 981 206 987
rect 266 981 324 987
rect -324 947 -312 981
rect -206 947 -194 981
rect -88 947 -76 981
rect 30 947 42 981
rect 148 947 160 981
rect 266 947 278 981
rect -324 941 -266 947
rect -206 941 -148 947
rect -88 941 -30 947
rect 30 941 88 947
rect 148 941 206 947
rect 266 941 324 947
rect -324 -947 -266 -941
rect -206 -947 -148 -941
rect -88 -947 -30 -941
rect 30 -947 88 -941
rect 148 -947 206 -941
rect 266 -947 324 -941
rect -324 -981 -312 -947
rect -206 -981 -194 -947
rect -88 -981 -76 -947
rect 30 -981 42 -947
rect 148 -981 160 -947
rect 266 -981 278 -947
rect -324 -987 -266 -981
rect -206 -987 -148 -981
rect -88 -987 -30 -981
rect 30 -987 88 -981
rect 148 -987 206 -981
rect 266 -987 324 -981
<< nwell >>
rect -521 -1119 521 1119
<< pmos >>
rect -325 -900 -265 900
rect -207 -900 -147 900
rect -89 -900 -29 900
rect 29 -900 89 900
rect 147 -900 207 900
rect 265 -900 325 900
<< pdiff >>
rect -383 888 -325 900
rect -383 -888 -371 888
rect -337 -888 -325 888
rect -383 -900 -325 -888
rect -265 888 -207 900
rect -265 -888 -253 888
rect -219 -888 -207 888
rect -265 -900 -207 -888
rect -147 888 -89 900
rect -147 -888 -135 888
rect -101 -888 -89 888
rect -147 -900 -89 -888
rect -29 888 29 900
rect -29 -888 -17 888
rect 17 -888 29 888
rect -29 -900 29 -888
rect 89 888 147 900
rect 89 -888 101 888
rect 135 -888 147 888
rect 89 -900 147 -888
rect 207 888 265 900
rect 207 -888 219 888
rect 253 -888 265 888
rect 207 -900 265 -888
rect 325 888 383 900
rect 325 -888 337 888
rect 371 -888 383 888
rect 325 -900 383 -888
<< pdiffc >>
rect -371 -888 -337 888
rect -253 -888 -219 888
rect -135 -888 -101 888
rect -17 -888 17 888
rect 101 -888 135 888
rect 219 -888 253 888
rect 337 -888 371 888
<< nsubdiff >>
rect -485 1049 -389 1083
rect 389 1049 485 1083
rect -485 987 -451 1049
rect 451 987 485 1049
rect -485 -1049 -451 -987
rect 451 -1049 485 -987
rect -485 -1083 -389 -1049
rect 389 -1083 485 -1049
<< nsubdiffcont >>
rect -389 1049 389 1083
rect -485 -987 -451 987
rect 451 -987 485 987
rect -389 -1083 389 -1049
<< poly >>
rect -328 981 -262 997
rect -328 947 -312 981
rect -278 947 -262 981
rect -328 931 -262 947
rect -210 981 -144 997
rect -210 947 -194 981
rect -160 947 -144 981
rect -210 931 -144 947
rect -92 981 -26 997
rect -92 947 -76 981
rect -42 947 -26 981
rect -92 931 -26 947
rect 26 981 92 997
rect 26 947 42 981
rect 76 947 92 981
rect 26 931 92 947
rect 144 981 210 997
rect 144 947 160 981
rect 194 947 210 981
rect 144 931 210 947
rect 262 981 328 997
rect 262 947 278 981
rect 312 947 328 981
rect 262 931 328 947
rect -325 900 -265 931
rect -207 900 -147 931
rect -89 900 -29 931
rect 29 900 89 931
rect 147 900 207 931
rect 265 900 325 931
rect -325 -931 -265 -900
rect -207 -931 -147 -900
rect -89 -931 -29 -900
rect 29 -931 89 -900
rect 147 -931 207 -900
rect 265 -931 325 -900
rect -328 -947 -262 -931
rect -328 -981 -312 -947
rect -278 -981 -262 -947
rect -328 -997 -262 -981
rect -210 -947 -144 -931
rect -210 -981 -194 -947
rect -160 -981 -144 -947
rect -210 -997 -144 -981
rect -92 -947 -26 -931
rect -92 -981 -76 -947
rect -42 -981 -26 -947
rect -92 -997 -26 -981
rect 26 -947 92 -931
rect 26 -981 42 -947
rect 76 -981 92 -947
rect 26 -997 92 -981
rect 144 -947 210 -931
rect 144 -981 160 -947
rect 194 -981 210 -947
rect 144 -997 210 -981
rect 262 -947 328 -931
rect 262 -981 278 -947
rect 312 -981 328 -947
rect 262 -997 328 -981
<< polycont >>
rect -312 947 -278 981
rect -194 947 -160 981
rect -76 947 -42 981
rect 42 947 76 981
rect 160 947 194 981
rect 278 947 312 981
rect -312 -981 -278 -947
rect -194 -981 -160 -947
rect -76 -981 -42 -947
rect 42 -981 76 -947
rect 160 -981 194 -947
rect 278 -981 312 -947
<< locali >>
rect -485 1049 -389 1083
rect 389 1049 485 1083
rect -485 987 -451 1049
rect 451 987 485 1049
rect -328 947 -312 981
rect -278 947 -262 981
rect -210 947 -194 981
rect -160 947 -144 981
rect -92 947 -76 981
rect -42 947 -26 981
rect 26 947 42 981
rect 76 947 92 981
rect 144 947 160 981
rect 194 947 210 981
rect 262 947 278 981
rect 312 947 328 981
rect -371 888 -337 904
rect -371 -904 -337 -888
rect -253 888 -219 904
rect -253 -904 -219 -888
rect -135 888 -101 904
rect -135 -904 -101 -888
rect -17 888 17 904
rect -17 -904 17 -888
rect 101 888 135 904
rect 101 -904 135 -888
rect 219 888 253 904
rect 219 -904 253 -888
rect 337 888 371 904
rect 337 -904 371 -888
rect -328 -981 -312 -947
rect -278 -981 -262 -947
rect -210 -981 -194 -947
rect -160 -981 -144 -947
rect -92 -981 -76 -947
rect -42 -981 -26 -947
rect 26 -981 42 -947
rect 76 -981 92 -947
rect 144 -981 160 -947
rect 194 -981 210 -947
rect 262 -981 278 -947
rect 312 -981 328 -947
rect -485 -1049 -451 -987
rect 451 -1049 485 -987
rect -485 -1083 -389 -1049
rect 389 -1083 485 -1049
<< viali >>
rect -312 947 -278 981
rect -194 947 -160 981
rect -76 947 -42 981
rect 42 947 76 981
rect 160 947 194 981
rect 278 947 312 981
rect -371 -888 -337 888
rect -253 -888 -219 888
rect -135 -888 -101 888
rect -17 -888 17 888
rect 101 -888 135 888
rect 219 -888 253 888
rect 337 -888 371 888
rect -312 -981 -278 -947
rect -194 -981 -160 -947
rect -76 -981 -42 -947
rect 42 -981 76 -947
rect 160 -981 194 -947
rect 278 -981 312 -947
<< metal1 >>
rect -324 981 -266 987
rect -324 947 -312 981
rect -278 947 -266 981
rect -324 941 -266 947
rect -206 981 -148 987
rect -206 947 -194 981
rect -160 947 -148 981
rect -206 941 -148 947
rect -88 981 -30 987
rect -88 947 -76 981
rect -42 947 -30 981
rect -88 941 -30 947
rect 30 981 88 987
rect 30 947 42 981
rect 76 947 88 981
rect 30 941 88 947
rect 148 981 206 987
rect 148 947 160 981
rect 194 947 206 981
rect 148 941 206 947
rect 266 981 324 987
rect 266 947 278 981
rect 312 947 324 981
rect 266 941 324 947
rect -377 888 -331 900
rect -377 -888 -371 888
rect -337 -888 -331 888
rect -377 -900 -331 -888
rect -259 888 -213 900
rect -259 -888 -253 888
rect -219 -888 -213 888
rect -259 -900 -213 -888
rect -141 888 -95 900
rect -141 -888 -135 888
rect -101 -888 -95 888
rect -141 -900 -95 -888
rect -23 888 23 900
rect -23 -888 -17 888
rect 17 -888 23 888
rect -23 -900 23 -888
rect 95 888 141 900
rect 95 -888 101 888
rect 135 -888 141 888
rect 95 -900 141 -888
rect 213 888 259 900
rect 213 -888 219 888
rect 253 -888 259 888
rect 213 -900 259 -888
rect 331 888 377 900
rect 331 -888 337 888
rect 371 -888 377 888
rect 331 -900 377 -888
rect -324 -947 -266 -941
rect -324 -981 -312 -947
rect -278 -981 -266 -947
rect -324 -987 -266 -981
rect -206 -947 -148 -941
rect -206 -981 -194 -947
rect -160 -981 -148 -947
rect -206 -987 -148 -981
rect -88 -947 -30 -941
rect -88 -981 -76 -947
rect -42 -981 -30 -947
rect -88 -987 -30 -981
rect 30 -947 88 -941
rect 30 -981 42 -947
rect 76 -981 88 -947
rect 30 -987 88 -981
rect 148 -947 206 -941
rect 148 -981 160 -947
rect 194 -981 206 -947
rect 148 -987 206 -981
rect 266 -947 324 -941
rect 266 -981 278 -947
rect 312 -981 324 -947
rect 266 -987 324 -981
<< properties >>
string FIXED_BBOX -468 -1066 468 1066
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 9 l 0.3 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
