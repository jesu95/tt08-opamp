magic
tech sky130A
magscale 1 2
timestamp 1723380300
<< nwell >>
rect -9067 -2737 9067 2737
<< pmos >>
rect -8871 118 -8751 2518
rect -8693 118 -8573 2518
rect -8515 118 -8395 2518
rect -8337 118 -8217 2518
rect -8159 118 -8039 2518
rect -7981 118 -7861 2518
rect -7803 118 -7683 2518
rect -7625 118 -7505 2518
rect -7447 118 -7327 2518
rect -7269 118 -7149 2518
rect -7091 118 -6971 2518
rect -6913 118 -6793 2518
rect -6735 118 -6615 2518
rect -6557 118 -6437 2518
rect -6379 118 -6259 2518
rect -6201 118 -6081 2518
rect -6023 118 -5903 2518
rect -5845 118 -5725 2518
rect -5667 118 -5547 2518
rect -5489 118 -5369 2518
rect -5311 118 -5191 2518
rect -5133 118 -5013 2518
rect -4955 118 -4835 2518
rect -4777 118 -4657 2518
rect -4599 118 -4479 2518
rect -4421 118 -4301 2518
rect -4243 118 -4123 2518
rect -4065 118 -3945 2518
rect -3887 118 -3767 2518
rect -3709 118 -3589 2518
rect -3531 118 -3411 2518
rect -3353 118 -3233 2518
rect -3175 118 -3055 2518
rect -2997 118 -2877 2518
rect -2819 118 -2699 2518
rect -2641 118 -2521 2518
rect -2463 118 -2343 2518
rect -2285 118 -2165 2518
rect -2107 118 -1987 2518
rect -1929 118 -1809 2518
rect -1751 118 -1631 2518
rect -1573 118 -1453 2518
rect -1395 118 -1275 2518
rect -1217 118 -1097 2518
rect -1039 118 -919 2518
rect -861 118 -741 2518
rect -683 118 -563 2518
rect -505 118 -385 2518
rect -327 118 -207 2518
rect -149 118 -29 2518
rect 29 118 149 2518
rect 207 118 327 2518
rect 385 118 505 2518
rect 563 118 683 2518
rect 741 118 861 2518
rect 919 118 1039 2518
rect 1097 118 1217 2518
rect 1275 118 1395 2518
rect 1453 118 1573 2518
rect 1631 118 1751 2518
rect 1809 118 1929 2518
rect 1987 118 2107 2518
rect 2165 118 2285 2518
rect 2343 118 2463 2518
rect 2521 118 2641 2518
rect 2699 118 2819 2518
rect 2877 118 2997 2518
rect 3055 118 3175 2518
rect 3233 118 3353 2518
rect 3411 118 3531 2518
rect 3589 118 3709 2518
rect 3767 118 3887 2518
rect 3945 118 4065 2518
rect 4123 118 4243 2518
rect 4301 118 4421 2518
rect 4479 118 4599 2518
rect 4657 118 4777 2518
rect 4835 118 4955 2518
rect 5013 118 5133 2518
rect 5191 118 5311 2518
rect 5369 118 5489 2518
rect 5547 118 5667 2518
rect 5725 118 5845 2518
rect 5903 118 6023 2518
rect 6081 118 6201 2518
rect 6259 118 6379 2518
rect 6437 118 6557 2518
rect 6615 118 6735 2518
rect 6793 118 6913 2518
rect 6971 118 7091 2518
rect 7149 118 7269 2518
rect 7327 118 7447 2518
rect 7505 118 7625 2518
rect 7683 118 7803 2518
rect 7861 118 7981 2518
rect 8039 118 8159 2518
rect 8217 118 8337 2518
rect 8395 118 8515 2518
rect 8573 118 8693 2518
rect 8751 118 8871 2518
rect -8871 -2518 -8751 -118
rect -8693 -2518 -8573 -118
rect -8515 -2518 -8395 -118
rect -8337 -2518 -8217 -118
rect -8159 -2518 -8039 -118
rect -7981 -2518 -7861 -118
rect -7803 -2518 -7683 -118
rect -7625 -2518 -7505 -118
rect -7447 -2518 -7327 -118
rect -7269 -2518 -7149 -118
rect -7091 -2518 -6971 -118
rect -6913 -2518 -6793 -118
rect -6735 -2518 -6615 -118
rect -6557 -2518 -6437 -118
rect -6379 -2518 -6259 -118
rect -6201 -2518 -6081 -118
rect -6023 -2518 -5903 -118
rect -5845 -2518 -5725 -118
rect -5667 -2518 -5547 -118
rect -5489 -2518 -5369 -118
rect -5311 -2518 -5191 -118
rect -5133 -2518 -5013 -118
rect -4955 -2518 -4835 -118
rect -4777 -2518 -4657 -118
rect -4599 -2518 -4479 -118
rect -4421 -2518 -4301 -118
rect -4243 -2518 -4123 -118
rect -4065 -2518 -3945 -118
rect -3887 -2518 -3767 -118
rect -3709 -2518 -3589 -118
rect -3531 -2518 -3411 -118
rect -3353 -2518 -3233 -118
rect -3175 -2518 -3055 -118
rect -2997 -2518 -2877 -118
rect -2819 -2518 -2699 -118
rect -2641 -2518 -2521 -118
rect -2463 -2518 -2343 -118
rect -2285 -2518 -2165 -118
rect -2107 -2518 -1987 -118
rect -1929 -2518 -1809 -118
rect -1751 -2518 -1631 -118
rect -1573 -2518 -1453 -118
rect -1395 -2518 -1275 -118
rect -1217 -2518 -1097 -118
rect -1039 -2518 -919 -118
rect -861 -2518 -741 -118
rect -683 -2518 -563 -118
rect -505 -2518 -385 -118
rect -327 -2518 -207 -118
rect -149 -2518 -29 -118
rect 29 -2518 149 -118
rect 207 -2518 327 -118
rect 385 -2518 505 -118
rect 563 -2518 683 -118
rect 741 -2518 861 -118
rect 919 -2518 1039 -118
rect 1097 -2518 1217 -118
rect 1275 -2518 1395 -118
rect 1453 -2518 1573 -118
rect 1631 -2518 1751 -118
rect 1809 -2518 1929 -118
rect 1987 -2518 2107 -118
rect 2165 -2518 2285 -118
rect 2343 -2518 2463 -118
rect 2521 -2518 2641 -118
rect 2699 -2518 2819 -118
rect 2877 -2518 2997 -118
rect 3055 -2518 3175 -118
rect 3233 -2518 3353 -118
rect 3411 -2518 3531 -118
rect 3589 -2518 3709 -118
rect 3767 -2518 3887 -118
rect 3945 -2518 4065 -118
rect 4123 -2518 4243 -118
rect 4301 -2518 4421 -118
rect 4479 -2518 4599 -118
rect 4657 -2518 4777 -118
rect 4835 -2518 4955 -118
rect 5013 -2518 5133 -118
rect 5191 -2518 5311 -118
rect 5369 -2518 5489 -118
rect 5547 -2518 5667 -118
rect 5725 -2518 5845 -118
rect 5903 -2518 6023 -118
rect 6081 -2518 6201 -118
rect 6259 -2518 6379 -118
rect 6437 -2518 6557 -118
rect 6615 -2518 6735 -118
rect 6793 -2518 6913 -118
rect 6971 -2518 7091 -118
rect 7149 -2518 7269 -118
rect 7327 -2518 7447 -118
rect 7505 -2518 7625 -118
rect 7683 -2518 7803 -118
rect 7861 -2518 7981 -118
rect 8039 -2518 8159 -118
rect 8217 -2518 8337 -118
rect 8395 -2518 8515 -118
rect 8573 -2518 8693 -118
rect 8751 -2518 8871 -118
<< pdiff >>
rect -8929 2506 -8871 2518
rect -8929 130 -8917 2506
rect -8883 130 -8871 2506
rect -8929 118 -8871 130
rect -8751 2506 -8693 2518
rect -8751 130 -8739 2506
rect -8705 130 -8693 2506
rect -8751 118 -8693 130
rect -8573 2506 -8515 2518
rect -8573 130 -8561 2506
rect -8527 130 -8515 2506
rect -8573 118 -8515 130
rect -8395 2506 -8337 2518
rect -8395 130 -8383 2506
rect -8349 130 -8337 2506
rect -8395 118 -8337 130
rect -8217 2506 -8159 2518
rect -8217 130 -8205 2506
rect -8171 130 -8159 2506
rect -8217 118 -8159 130
rect -8039 2506 -7981 2518
rect -8039 130 -8027 2506
rect -7993 130 -7981 2506
rect -8039 118 -7981 130
rect -7861 2506 -7803 2518
rect -7861 130 -7849 2506
rect -7815 130 -7803 2506
rect -7861 118 -7803 130
rect -7683 2506 -7625 2518
rect -7683 130 -7671 2506
rect -7637 130 -7625 2506
rect -7683 118 -7625 130
rect -7505 2506 -7447 2518
rect -7505 130 -7493 2506
rect -7459 130 -7447 2506
rect -7505 118 -7447 130
rect -7327 2506 -7269 2518
rect -7327 130 -7315 2506
rect -7281 130 -7269 2506
rect -7327 118 -7269 130
rect -7149 2506 -7091 2518
rect -7149 130 -7137 2506
rect -7103 130 -7091 2506
rect -7149 118 -7091 130
rect -6971 2506 -6913 2518
rect -6971 130 -6959 2506
rect -6925 130 -6913 2506
rect -6971 118 -6913 130
rect -6793 2506 -6735 2518
rect -6793 130 -6781 2506
rect -6747 130 -6735 2506
rect -6793 118 -6735 130
rect -6615 2506 -6557 2518
rect -6615 130 -6603 2506
rect -6569 130 -6557 2506
rect -6615 118 -6557 130
rect -6437 2506 -6379 2518
rect -6437 130 -6425 2506
rect -6391 130 -6379 2506
rect -6437 118 -6379 130
rect -6259 2506 -6201 2518
rect -6259 130 -6247 2506
rect -6213 130 -6201 2506
rect -6259 118 -6201 130
rect -6081 2506 -6023 2518
rect -6081 130 -6069 2506
rect -6035 130 -6023 2506
rect -6081 118 -6023 130
rect -5903 2506 -5845 2518
rect -5903 130 -5891 2506
rect -5857 130 -5845 2506
rect -5903 118 -5845 130
rect -5725 2506 -5667 2518
rect -5725 130 -5713 2506
rect -5679 130 -5667 2506
rect -5725 118 -5667 130
rect -5547 2506 -5489 2518
rect -5547 130 -5535 2506
rect -5501 130 -5489 2506
rect -5547 118 -5489 130
rect -5369 2506 -5311 2518
rect -5369 130 -5357 2506
rect -5323 130 -5311 2506
rect -5369 118 -5311 130
rect -5191 2506 -5133 2518
rect -5191 130 -5179 2506
rect -5145 130 -5133 2506
rect -5191 118 -5133 130
rect -5013 2506 -4955 2518
rect -5013 130 -5001 2506
rect -4967 130 -4955 2506
rect -5013 118 -4955 130
rect -4835 2506 -4777 2518
rect -4835 130 -4823 2506
rect -4789 130 -4777 2506
rect -4835 118 -4777 130
rect -4657 2506 -4599 2518
rect -4657 130 -4645 2506
rect -4611 130 -4599 2506
rect -4657 118 -4599 130
rect -4479 2506 -4421 2518
rect -4479 130 -4467 2506
rect -4433 130 -4421 2506
rect -4479 118 -4421 130
rect -4301 2506 -4243 2518
rect -4301 130 -4289 2506
rect -4255 130 -4243 2506
rect -4301 118 -4243 130
rect -4123 2506 -4065 2518
rect -4123 130 -4111 2506
rect -4077 130 -4065 2506
rect -4123 118 -4065 130
rect -3945 2506 -3887 2518
rect -3945 130 -3933 2506
rect -3899 130 -3887 2506
rect -3945 118 -3887 130
rect -3767 2506 -3709 2518
rect -3767 130 -3755 2506
rect -3721 130 -3709 2506
rect -3767 118 -3709 130
rect -3589 2506 -3531 2518
rect -3589 130 -3577 2506
rect -3543 130 -3531 2506
rect -3589 118 -3531 130
rect -3411 2506 -3353 2518
rect -3411 130 -3399 2506
rect -3365 130 -3353 2506
rect -3411 118 -3353 130
rect -3233 2506 -3175 2518
rect -3233 130 -3221 2506
rect -3187 130 -3175 2506
rect -3233 118 -3175 130
rect -3055 2506 -2997 2518
rect -3055 130 -3043 2506
rect -3009 130 -2997 2506
rect -3055 118 -2997 130
rect -2877 2506 -2819 2518
rect -2877 130 -2865 2506
rect -2831 130 -2819 2506
rect -2877 118 -2819 130
rect -2699 2506 -2641 2518
rect -2699 130 -2687 2506
rect -2653 130 -2641 2506
rect -2699 118 -2641 130
rect -2521 2506 -2463 2518
rect -2521 130 -2509 2506
rect -2475 130 -2463 2506
rect -2521 118 -2463 130
rect -2343 2506 -2285 2518
rect -2343 130 -2331 2506
rect -2297 130 -2285 2506
rect -2343 118 -2285 130
rect -2165 2506 -2107 2518
rect -2165 130 -2153 2506
rect -2119 130 -2107 2506
rect -2165 118 -2107 130
rect -1987 2506 -1929 2518
rect -1987 130 -1975 2506
rect -1941 130 -1929 2506
rect -1987 118 -1929 130
rect -1809 2506 -1751 2518
rect -1809 130 -1797 2506
rect -1763 130 -1751 2506
rect -1809 118 -1751 130
rect -1631 2506 -1573 2518
rect -1631 130 -1619 2506
rect -1585 130 -1573 2506
rect -1631 118 -1573 130
rect -1453 2506 -1395 2518
rect -1453 130 -1441 2506
rect -1407 130 -1395 2506
rect -1453 118 -1395 130
rect -1275 2506 -1217 2518
rect -1275 130 -1263 2506
rect -1229 130 -1217 2506
rect -1275 118 -1217 130
rect -1097 2506 -1039 2518
rect -1097 130 -1085 2506
rect -1051 130 -1039 2506
rect -1097 118 -1039 130
rect -919 2506 -861 2518
rect -919 130 -907 2506
rect -873 130 -861 2506
rect -919 118 -861 130
rect -741 2506 -683 2518
rect -741 130 -729 2506
rect -695 130 -683 2506
rect -741 118 -683 130
rect -563 2506 -505 2518
rect -563 130 -551 2506
rect -517 130 -505 2506
rect -563 118 -505 130
rect -385 2506 -327 2518
rect -385 130 -373 2506
rect -339 130 -327 2506
rect -385 118 -327 130
rect -207 2506 -149 2518
rect -207 130 -195 2506
rect -161 130 -149 2506
rect -207 118 -149 130
rect -29 2506 29 2518
rect -29 130 -17 2506
rect 17 130 29 2506
rect -29 118 29 130
rect 149 2506 207 2518
rect 149 130 161 2506
rect 195 130 207 2506
rect 149 118 207 130
rect 327 2506 385 2518
rect 327 130 339 2506
rect 373 130 385 2506
rect 327 118 385 130
rect 505 2506 563 2518
rect 505 130 517 2506
rect 551 130 563 2506
rect 505 118 563 130
rect 683 2506 741 2518
rect 683 130 695 2506
rect 729 130 741 2506
rect 683 118 741 130
rect 861 2506 919 2518
rect 861 130 873 2506
rect 907 130 919 2506
rect 861 118 919 130
rect 1039 2506 1097 2518
rect 1039 130 1051 2506
rect 1085 130 1097 2506
rect 1039 118 1097 130
rect 1217 2506 1275 2518
rect 1217 130 1229 2506
rect 1263 130 1275 2506
rect 1217 118 1275 130
rect 1395 2506 1453 2518
rect 1395 130 1407 2506
rect 1441 130 1453 2506
rect 1395 118 1453 130
rect 1573 2506 1631 2518
rect 1573 130 1585 2506
rect 1619 130 1631 2506
rect 1573 118 1631 130
rect 1751 2506 1809 2518
rect 1751 130 1763 2506
rect 1797 130 1809 2506
rect 1751 118 1809 130
rect 1929 2506 1987 2518
rect 1929 130 1941 2506
rect 1975 130 1987 2506
rect 1929 118 1987 130
rect 2107 2506 2165 2518
rect 2107 130 2119 2506
rect 2153 130 2165 2506
rect 2107 118 2165 130
rect 2285 2506 2343 2518
rect 2285 130 2297 2506
rect 2331 130 2343 2506
rect 2285 118 2343 130
rect 2463 2506 2521 2518
rect 2463 130 2475 2506
rect 2509 130 2521 2506
rect 2463 118 2521 130
rect 2641 2506 2699 2518
rect 2641 130 2653 2506
rect 2687 130 2699 2506
rect 2641 118 2699 130
rect 2819 2506 2877 2518
rect 2819 130 2831 2506
rect 2865 130 2877 2506
rect 2819 118 2877 130
rect 2997 2506 3055 2518
rect 2997 130 3009 2506
rect 3043 130 3055 2506
rect 2997 118 3055 130
rect 3175 2506 3233 2518
rect 3175 130 3187 2506
rect 3221 130 3233 2506
rect 3175 118 3233 130
rect 3353 2506 3411 2518
rect 3353 130 3365 2506
rect 3399 130 3411 2506
rect 3353 118 3411 130
rect 3531 2506 3589 2518
rect 3531 130 3543 2506
rect 3577 130 3589 2506
rect 3531 118 3589 130
rect 3709 2506 3767 2518
rect 3709 130 3721 2506
rect 3755 130 3767 2506
rect 3709 118 3767 130
rect 3887 2506 3945 2518
rect 3887 130 3899 2506
rect 3933 130 3945 2506
rect 3887 118 3945 130
rect 4065 2506 4123 2518
rect 4065 130 4077 2506
rect 4111 130 4123 2506
rect 4065 118 4123 130
rect 4243 2506 4301 2518
rect 4243 130 4255 2506
rect 4289 130 4301 2506
rect 4243 118 4301 130
rect 4421 2506 4479 2518
rect 4421 130 4433 2506
rect 4467 130 4479 2506
rect 4421 118 4479 130
rect 4599 2506 4657 2518
rect 4599 130 4611 2506
rect 4645 130 4657 2506
rect 4599 118 4657 130
rect 4777 2506 4835 2518
rect 4777 130 4789 2506
rect 4823 130 4835 2506
rect 4777 118 4835 130
rect 4955 2506 5013 2518
rect 4955 130 4967 2506
rect 5001 130 5013 2506
rect 4955 118 5013 130
rect 5133 2506 5191 2518
rect 5133 130 5145 2506
rect 5179 130 5191 2506
rect 5133 118 5191 130
rect 5311 2506 5369 2518
rect 5311 130 5323 2506
rect 5357 130 5369 2506
rect 5311 118 5369 130
rect 5489 2506 5547 2518
rect 5489 130 5501 2506
rect 5535 130 5547 2506
rect 5489 118 5547 130
rect 5667 2506 5725 2518
rect 5667 130 5679 2506
rect 5713 130 5725 2506
rect 5667 118 5725 130
rect 5845 2506 5903 2518
rect 5845 130 5857 2506
rect 5891 130 5903 2506
rect 5845 118 5903 130
rect 6023 2506 6081 2518
rect 6023 130 6035 2506
rect 6069 130 6081 2506
rect 6023 118 6081 130
rect 6201 2506 6259 2518
rect 6201 130 6213 2506
rect 6247 130 6259 2506
rect 6201 118 6259 130
rect 6379 2506 6437 2518
rect 6379 130 6391 2506
rect 6425 130 6437 2506
rect 6379 118 6437 130
rect 6557 2506 6615 2518
rect 6557 130 6569 2506
rect 6603 130 6615 2506
rect 6557 118 6615 130
rect 6735 2506 6793 2518
rect 6735 130 6747 2506
rect 6781 130 6793 2506
rect 6735 118 6793 130
rect 6913 2506 6971 2518
rect 6913 130 6925 2506
rect 6959 130 6971 2506
rect 6913 118 6971 130
rect 7091 2506 7149 2518
rect 7091 130 7103 2506
rect 7137 130 7149 2506
rect 7091 118 7149 130
rect 7269 2506 7327 2518
rect 7269 130 7281 2506
rect 7315 130 7327 2506
rect 7269 118 7327 130
rect 7447 2506 7505 2518
rect 7447 130 7459 2506
rect 7493 130 7505 2506
rect 7447 118 7505 130
rect 7625 2506 7683 2518
rect 7625 130 7637 2506
rect 7671 130 7683 2506
rect 7625 118 7683 130
rect 7803 2506 7861 2518
rect 7803 130 7815 2506
rect 7849 130 7861 2506
rect 7803 118 7861 130
rect 7981 2506 8039 2518
rect 7981 130 7993 2506
rect 8027 130 8039 2506
rect 7981 118 8039 130
rect 8159 2506 8217 2518
rect 8159 130 8171 2506
rect 8205 130 8217 2506
rect 8159 118 8217 130
rect 8337 2506 8395 2518
rect 8337 130 8349 2506
rect 8383 130 8395 2506
rect 8337 118 8395 130
rect 8515 2506 8573 2518
rect 8515 130 8527 2506
rect 8561 130 8573 2506
rect 8515 118 8573 130
rect 8693 2506 8751 2518
rect 8693 130 8705 2506
rect 8739 130 8751 2506
rect 8693 118 8751 130
rect 8871 2506 8929 2518
rect 8871 130 8883 2506
rect 8917 130 8929 2506
rect 8871 118 8929 130
rect -8929 -130 -8871 -118
rect -8929 -2506 -8917 -130
rect -8883 -2506 -8871 -130
rect -8929 -2518 -8871 -2506
rect -8751 -130 -8693 -118
rect -8751 -2506 -8739 -130
rect -8705 -2506 -8693 -130
rect -8751 -2518 -8693 -2506
rect -8573 -130 -8515 -118
rect -8573 -2506 -8561 -130
rect -8527 -2506 -8515 -130
rect -8573 -2518 -8515 -2506
rect -8395 -130 -8337 -118
rect -8395 -2506 -8383 -130
rect -8349 -2506 -8337 -130
rect -8395 -2518 -8337 -2506
rect -8217 -130 -8159 -118
rect -8217 -2506 -8205 -130
rect -8171 -2506 -8159 -130
rect -8217 -2518 -8159 -2506
rect -8039 -130 -7981 -118
rect -8039 -2506 -8027 -130
rect -7993 -2506 -7981 -130
rect -8039 -2518 -7981 -2506
rect -7861 -130 -7803 -118
rect -7861 -2506 -7849 -130
rect -7815 -2506 -7803 -130
rect -7861 -2518 -7803 -2506
rect -7683 -130 -7625 -118
rect -7683 -2506 -7671 -130
rect -7637 -2506 -7625 -130
rect -7683 -2518 -7625 -2506
rect -7505 -130 -7447 -118
rect -7505 -2506 -7493 -130
rect -7459 -2506 -7447 -130
rect -7505 -2518 -7447 -2506
rect -7327 -130 -7269 -118
rect -7327 -2506 -7315 -130
rect -7281 -2506 -7269 -130
rect -7327 -2518 -7269 -2506
rect -7149 -130 -7091 -118
rect -7149 -2506 -7137 -130
rect -7103 -2506 -7091 -130
rect -7149 -2518 -7091 -2506
rect -6971 -130 -6913 -118
rect -6971 -2506 -6959 -130
rect -6925 -2506 -6913 -130
rect -6971 -2518 -6913 -2506
rect -6793 -130 -6735 -118
rect -6793 -2506 -6781 -130
rect -6747 -2506 -6735 -130
rect -6793 -2518 -6735 -2506
rect -6615 -130 -6557 -118
rect -6615 -2506 -6603 -130
rect -6569 -2506 -6557 -130
rect -6615 -2518 -6557 -2506
rect -6437 -130 -6379 -118
rect -6437 -2506 -6425 -130
rect -6391 -2506 -6379 -130
rect -6437 -2518 -6379 -2506
rect -6259 -130 -6201 -118
rect -6259 -2506 -6247 -130
rect -6213 -2506 -6201 -130
rect -6259 -2518 -6201 -2506
rect -6081 -130 -6023 -118
rect -6081 -2506 -6069 -130
rect -6035 -2506 -6023 -130
rect -6081 -2518 -6023 -2506
rect -5903 -130 -5845 -118
rect -5903 -2506 -5891 -130
rect -5857 -2506 -5845 -130
rect -5903 -2518 -5845 -2506
rect -5725 -130 -5667 -118
rect -5725 -2506 -5713 -130
rect -5679 -2506 -5667 -130
rect -5725 -2518 -5667 -2506
rect -5547 -130 -5489 -118
rect -5547 -2506 -5535 -130
rect -5501 -2506 -5489 -130
rect -5547 -2518 -5489 -2506
rect -5369 -130 -5311 -118
rect -5369 -2506 -5357 -130
rect -5323 -2506 -5311 -130
rect -5369 -2518 -5311 -2506
rect -5191 -130 -5133 -118
rect -5191 -2506 -5179 -130
rect -5145 -2506 -5133 -130
rect -5191 -2518 -5133 -2506
rect -5013 -130 -4955 -118
rect -5013 -2506 -5001 -130
rect -4967 -2506 -4955 -130
rect -5013 -2518 -4955 -2506
rect -4835 -130 -4777 -118
rect -4835 -2506 -4823 -130
rect -4789 -2506 -4777 -130
rect -4835 -2518 -4777 -2506
rect -4657 -130 -4599 -118
rect -4657 -2506 -4645 -130
rect -4611 -2506 -4599 -130
rect -4657 -2518 -4599 -2506
rect -4479 -130 -4421 -118
rect -4479 -2506 -4467 -130
rect -4433 -2506 -4421 -130
rect -4479 -2518 -4421 -2506
rect -4301 -130 -4243 -118
rect -4301 -2506 -4289 -130
rect -4255 -2506 -4243 -130
rect -4301 -2518 -4243 -2506
rect -4123 -130 -4065 -118
rect -4123 -2506 -4111 -130
rect -4077 -2506 -4065 -130
rect -4123 -2518 -4065 -2506
rect -3945 -130 -3887 -118
rect -3945 -2506 -3933 -130
rect -3899 -2506 -3887 -130
rect -3945 -2518 -3887 -2506
rect -3767 -130 -3709 -118
rect -3767 -2506 -3755 -130
rect -3721 -2506 -3709 -130
rect -3767 -2518 -3709 -2506
rect -3589 -130 -3531 -118
rect -3589 -2506 -3577 -130
rect -3543 -2506 -3531 -130
rect -3589 -2518 -3531 -2506
rect -3411 -130 -3353 -118
rect -3411 -2506 -3399 -130
rect -3365 -2506 -3353 -130
rect -3411 -2518 -3353 -2506
rect -3233 -130 -3175 -118
rect -3233 -2506 -3221 -130
rect -3187 -2506 -3175 -130
rect -3233 -2518 -3175 -2506
rect -3055 -130 -2997 -118
rect -3055 -2506 -3043 -130
rect -3009 -2506 -2997 -130
rect -3055 -2518 -2997 -2506
rect -2877 -130 -2819 -118
rect -2877 -2506 -2865 -130
rect -2831 -2506 -2819 -130
rect -2877 -2518 -2819 -2506
rect -2699 -130 -2641 -118
rect -2699 -2506 -2687 -130
rect -2653 -2506 -2641 -130
rect -2699 -2518 -2641 -2506
rect -2521 -130 -2463 -118
rect -2521 -2506 -2509 -130
rect -2475 -2506 -2463 -130
rect -2521 -2518 -2463 -2506
rect -2343 -130 -2285 -118
rect -2343 -2506 -2331 -130
rect -2297 -2506 -2285 -130
rect -2343 -2518 -2285 -2506
rect -2165 -130 -2107 -118
rect -2165 -2506 -2153 -130
rect -2119 -2506 -2107 -130
rect -2165 -2518 -2107 -2506
rect -1987 -130 -1929 -118
rect -1987 -2506 -1975 -130
rect -1941 -2506 -1929 -130
rect -1987 -2518 -1929 -2506
rect -1809 -130 -1751 -118
rect -1809 -2506 -1797 -130
rect -1763 -2506 -1751 -130
rect -1809 -2518 -1751 -2506
rect -1631 -130 -1573 -118
rect -1631 -2506 -1619 -130
rect -1585 -2506 -1573 -130
rect -1631 -2518 -1573 -2506
rect -1453 -130 -1395 -118
rect -1453 -2506 -1441 -130
rect -1407 -2506 -1395 -130
rect -1453 -2518 -1395 -2506
rect -1275 -130 -1217 -118
rect -1275 -2506 -1263 -130
rect -1229 -2506 -1217 -130
rect -1275 -2518 -1217 -2506
rect -1097 -130 -1039 -118
rect -1097 -2506 -1085 -130
rect -1051 -2506 -1039 -130
rect -1097 -2518 -1039 -2506
rect -919 -130 -861 -118
rect -919 -2506 -907 -130
rect -873 -2506 -861 -130
rect -919 -2518 -861 -2506
rect -741 -130 -683 -118
rect -741 -2506 -729 -130
rect -695 -2506 -683 -130
rect -741 -2518 -683 -2506
rect -563 -130 -505 -118
rect -563 -2506 -551 -130
rect -517 -2506 -505 -130
rect -563 -2518 -505 -2506
rect -385 -130 -327 -118
rect -385 -2506 -373 -130
rect -339 -2506 -327 -130
rect -385 -2518 -327 -2506
rect -207 -130 -149 -118
rect -207 -2506 -195 -130
rect -161 -2506 -149 -130
rect -207 -2518 -149 -2506
rect -29 -130 29 -118
rect -29 -2506 -17 -130
rect 17 -2506 29 -130
rect -29 -2518 29 -2506
rect 149 -130 207 -118
rect 149 -2506 161 -130
rect 195 -2506 207 -130
rect 149 -2518 207 -2506
rect 327 -130 385 -118
rect 327 -2506 339 -130
rect 373 -2506 385 -130
rect 327 -2518 385 -2506
rect 505 -130 563 -118
rect 505 -2506 517 -130
rect 551 -2506 563 -130
rect 505 -2518 563 -2506
rect 683 -130 741 -118
rect 683 -2506 695 -130
rect 729 -2506 741 -130
rect 683 -2518 741 -2506
rect 861 -130 919 -118
rect 861 -2506 873 -130
rect 907 -2506 919 -130
rect 861 -2518 919 -2506
rect 1039 -130 1097 -118
rect 1039 -2506 1051 -130
rect 1085 -2506 1097 -130
rect 1039 -2518 1097 -2506
rect 1217 -130 1275 -118
rect 1217 -2506 1229 -130
rect 1263 -2506 1275 -130
rect 1217 -2518 1275 -2506
rect 1395 -130 1453 -118
rect 1395 -2506 1407 -130
rect 1441 -2506 1453 -130
rect 1395 -2518 1453 -2506
rect 1573 -130 1631 -118
rect 1573 -2506 1585 -130
rect 1619 -2506 1631 -130
rect 1573 -2518 1631 -2506
rect 1751 -130 1809 -118
rect 1751 -2506 1763 -130
rect 1797 -2506 1809 -130
rect 1751 -2518 1809 -2506
rect 1929 -130 1987 -118
rect 1929 -2506 1941 -130
rect 1975 -2506 1987 -130
rect 1929 -2518 1987 -2506
rect 2107 -130 2165 -118
rect 2107 -2506 2119 -130
rect 2153 -2506 2165 -130
rect 2107 -2518 2165 -2506
rect 2285 -130 2343 -118
rect 2285 -2506 2297 -130
rect 2331 -2506 2343 -130
rect 2285 -2518 2343 -2506
rect 2463 -130 2521 -118
rect 2463 -2506 2475 -130
rect 2509 -2506 2521 -130
rect 2463 -2518 2521 -2506
rect 2641 -130 2699 -118
rect 2641 -2506 2653 -130
rect 2687 -2506 2699 -130
rect 2641 -2518 2699 -2506
rect 2819 -130 2877 -118
rect 2819 -2506 2831 -130
rect 2865 -2506 2877 -130
rect 2819 -2518 2877 -2506
rect 2997 -130 3055 -118
rect 2997 -2506 3009 -130
rect 3043 -2506 3055 -130
rect 2997 -2518 3055 -2506
rect 3175 -130 3233 -118
rect 3175 -2506 3187 -130
rect 3221 -2506 3233 -130
rect 3175 -2518 3233 -2506
rect 3353 -130 3411 -118
rect 3353 -2506 3365 -130
rect 3399 -2506 3411 -130
rect 3353 -2518 3411 -2506
rect 3531 -130 3589 -118
rect 3531 -2506 3543 -130
rect 3577 -2506 3589 -130
rect 3531 -2518 3589 -2506
rect 3709 -130 3767 -118
rect 3709 -2506 3721 -130
rect 3755 -2506 3767 -130
rect 3709 -2518 3767 -2506
rect 3887 -130 3945 -118
rect 3887 -2506 3899 -130
rect 3933 -2506 3945 -130
rect 3887 -2518 3945 -2506
rect 4065 -130 4123 -118
rect 4065 -2506 4077 -130
rect 4111 -2506 4123 -130
rect 4065 -2518 4123 -2506
rect 4243 -130 4301 -118
rect 4243 -2506 4255 -130
rect 4289 -2506 4301 -130
rect 4243 -2518 4301 -2506
rect 4421 -130 4479 -118
rect 4421 -2506 4433 -130
rect 4467 -2506 4479 -130
rect 4421 -2518 4479 -2506
rect 4599 -130 4657 -118
rect 4599 -2506 4611 -130
rect 4645 -2506 4657 -130
rect 4599 -2518 4657 -2506
rect 4777 -130 4835 -118
rect 4777 -2506 4789 -130
rect 4823 -2506 4835 -130
rect 4777 -2518 4835 -2506
rect 4955 -130 5013 -118
rect 4955 -2506 4967 -130
rect 5001 -2506 5013 -130
rect 4955 -2518 5013 -2506
rect 5133 -130 5191 -118
rect 5133 -2506 5145 -130
rect 5179 -2506 5191 -130
rect 5133 -2518 5191 -2506
rect 5311 -130 5369 -118
rect 5311 -2506 5323 -130
rect 5357 -2506 5369 -130
rect 5311 -2518 5369 -2506
rect 5489 -130 5547 -118
rect 5489 -2506 5501 -130
rect 5535 -2506 5547 -130
rect 5489 -2518 5547 -2506
rect 5667 -130 5725 -118
rect 5667 -2506 5679 -130
rect 5713 -2506 5725 -130
rect 5667 -2518 5725 -2506
rect 5845 -130 5903 -118
rect 5845 -2506 5857 -130
rect 5891 -2506 5903 -130
rect 5845 -2518 5903 -2506
rect 6023 -130 6081 -118
rect 6023 -2506 6035 -130
rect 6069 -2506 6081 -130
rect 6023 -2518 6081 -2506
rect 6201 -130 6259 -118
rect 6201 -2506 6213 -130
rect 6247 -2506 6259 -130
rect 6201 -2518 6259 -2506
rect 6379 -130 6437 -118
rect 6379 -2506 6391 -130
rect 6425 -2506 6437 -130
rect 6379 -2518 6437 -2506
rect 6557 -130 6615 -118
rect 6557 -2506 6569 -130
rect 6603 -2506 6615 -130
rect 6557 -2518 6615 -2506
rect 6735 -130 6793 -118
rect 6735 -2506 6747 -130
rect 6781 -2506 6793 -130
rect 6735 -2518 6793 -2506
rect 6913 -130 6971 -118
rect 6913 -2506 6925 -130
rect 6959 -2506 6971 -130
rect 6913 -2518 6971 -2506
rect 7091 -130 7149 -118
rect 7091 -2506 7103 -130
rect 7137 -2506 7149 -130
rect 7091 -2518 7149 -2506
rect 7269 -130 7327 -118
rect 7269 -2506 7281 -130
rect 7315 -2506 7327 -130
rect 7269 -2518 7327 -2506
rect 7447 -130 7505 -118
rect 7447 -2506 7459 -130
rect 7493 -2506 7505 -130
rect 7447 -2518 7505 -2506
rect 7625 -130 7683 -118
rect 7625 -2506 7637 -130
rect 7671 -2506 7683 -130
rect 7625 -2518 7683 -2506
rect 7803 -130 7861 -118
rect 7803 -2506 7815 -130
rect 7849 -2506 7861 -130
rect 7803 -2518 7861 -2506
rect 7981 -130 8039 -118
rect 7981 -2506 7993 -130
rect 8027 -2506 8039 -130
rect 7981 -2518 8039 -2506
rect 8159 -130 8217 -118
rect 8159 -2506 8171 -130
rect 8205 -2506 8217 -130
rect 8159 -2518 8217 -2506
rect 8337 -130 8395 -118
rect 8337 -2506 8349 -130
rect 8383 -2506 8395 -130
rect 8337 -2518 8395 -2506
rect 8515 -130 8573 -118
rect 8515 -2506 8527 -130
rect 8561 -2506 8573 -130
rect 8515 -2518 8573 -2506
rect 8693 -130 8751 -118
rect 8693 -2506 8705 -130
rect 8739 -2506 8751 -130
rect 8693 -2518 8751 -2506
rect 8871 -130 8929 -118
rect 8871 -2506 8883 -130
rect 8917 -2506 8929 -130
rect 8871 -2518 8929 -2506
<< pdiffc >>
rect -8917 130 -8883 2506
rect -8739 130 -8705 2506
rect -8561 130 -8527 2506
rect -8383 130 -8349 2506
rect -8205 130 -8171 2506
rect -8027 130 -7993 2506
rect -7849 130 -7815 2506
rect -7671 130 -7637 2506
rect -7493 130 -7459 2506
rect -7315 130 -7281 2506
rect -7137 130 -7103 2506
rect -6959 130 -6925 2506
rect -6781 130 -6747 2506
rect -6603 130 -6569 2506
rect -6425 130 -6391 2506
rect -6247 130 -6213 2506
rect -6069 130 -6035 2506
rect -5891 130 -5857 2506
rect -5713 130 -5679 2506
rect -5535 130 -5501 2506
rect -5357 130 -5323 2506
rect -5179 130 -5145 2506
rect -5001 130 -4967 2506
rect -4823 130 -4789 2506
rect -4645 130 -4611 2506
rect -4467 130 -4433 2506
rect -4289 130 -4255 2506
rect -4111 130 -4077 2506
rect -3933 130 -3899 2506
rect -3755 130 -3721 2506
rect -3577 130 -3543 2506
rect -3399 130 -3365 2506
rect -3221 130 -3187 2506
rect -3043 130 -3009 2506
rect -2865 130 -2831 2506
rect -2687 130 -2653 2506
rect -2509 130 -2475 2506
rect -2331 130 -2297 2506
rect -2153 130 -2119 2506
rect -1975 130 -1941 2506
rect -1797 130 -1763 2506
rect -1619 130 -1585 2506
rect -1441 130 -1407 2506
rect -1263 130 -1229 2506
rect -1085 130 -1051 2506
rect -907 130 -873 2506
rect -729 130 -695 2506
rect -551 130 -517 2506
rect -373 130 -339 2506
rect -195 130 -161 2506
rect -17 130 17 2506
rect 161 130 195 2506
rect 339 130 373 2506
rect 517 130 551 2506
rect 695 130 729 2506
rect 873 130 907 2506
rect 1051 130 1085 2506
rect 1229 130 1263 2506
rect 1407 130 1441 2506
rect 1585 130 1619 2506
rect 1763 130 1797 2506
rect 1941 130 1975 2506
rect 2119 130 2153 2506
rect 2297 130 2331 2506
rect 2475 130 2509 2506
rect 2653 130 2687 2506
rect 2831 130 2865 2506
rect 3009 130 3043 2506
rect 3187 130 3221 2506
rect 3365 130 3399 2506
rect 3543 130 3577 2506
rect 3721 130 3755 2506
rect 3899 130 3933 2506
rect 4077 130 4111 2506
rect 4255 130 4289 2506
rect 4433 130 4467 2506
rect 4611 130 4645 2506
rect 4789 130 4823 2506
rect 4967 130 5001 2506
rect 5145 130 5179 2506
rect 5323 130 5357 2506
rect 5501 130 5535 2506
rect 5679 130 5713 2506
rect 5857 130 5891 2506
rect 6035 130 6069 2506
rect 6213 130 6247 2506
rect 6391 130 6425 2506
rect 6569 130 6603 2506
rect 6747 130 6781 2506
rect 6925 130 6959 2506
rect 7103 130 7137 2506
rect 7281 130 7315 2506
rect 7459 130 7493 2506
rect 7637 130 7671 2506
rect 7815 130 7849 2506
rect 7993 130 8027 2506
rect 8171 130 8205 2506
rect 8349 130 8383 2506
rect 8527 130 8561 2506
rect 8705 130 8739 2506
rect 8883 130 8917 2506
rect -8917 -2506 -8883 -130
rect -8739 -2506 -8705 -130
rect -8561 -2506 -8527 -130
rect -8383 -2506 -8349 -130
rect -8205 -2506 -8171 -130
rect -8027 -2506 -7993 -130
rect -7849 -2506 -7815 -130
rect -7671 -2506 -7637 -130
rect -7493 -2506 -7459 -130
rect -7315 -2506 -7281 -130
rect -7137 -2506 -7103 -130
rect -6959 -2506 -6925 -130
rect -6781 -2506 -6747 -130
rect -6603 -2506 -6569 -130
rect -6425 -2506 -6391 -130
rect -6247 -2506 -6213 -130
rect -6069 -2506 -6035 -130
rect -5891 -2506 -5857 -130
rect -5713 -2506 -5679 -130
rect -5535 -2506 -5501 -130
rect -5357 -2506 -5323 -130
rect -5179 -2506 -5145 -130
rect -5001 -2506 -4967 -130
rect -4823 -2506 -4789 -130
rect -4645 -2506 -4611 -130
rect -4467 -2506 -4433 -130
rect -4289 -2506 -4255 -130
rect -4111 -2506 -4077 -130
rect -3933 -2506 -3899 -130
rect -3755 -2506 -3721 -130
rect -3577 -2506 -3543 -130
rect -3399 -2506 -3365 -130
rect -3221 -2506 -3187 -130
rect -3043 -2506 -3009 -130
rect -2865 -2506 -2831 -130
rect -2687 -2506 -2653 -130
rect -2509 -2506 -2475 -130
rect -2331 -2506 -2297 -130
rect -2153 -2506 -2119 -130
rect -1975 -2506 -1941 -130
rect -1797 -2506 -1763 -130
rect -1619 -2506 -1585 -130
rect -1441 -2506 -1407 -130
rect -1263 -2506 -1229 -130
rect -1085 -2506 -1051 -130
rect -907 -2506 -873 -130
rect -729 -2506 -695 -130
rect -551 -2506 -517 -130
rect -373 -2506 -339 -130
rect -195 -2506 -161 -130
rect -17 -2506 17 -130
rect 161 -2506 195 -130
rect 339 -2506 373 -130
rect 517 -2506 551 -130
rect 695 -2506 729 -130
rect 873 -2506 907 -130
rect 1051 -2506 1085 -130
rect 1229 -2506 1263 -130
rect 1407 -2506 1441 -130
rect 1585 -2506 1619 -130
rect 1763 -2506 1797 -130
rect 1941 -2506 1975 -130
rect 2119 -2506 2153 -130
rect 2297 -2506 2331 -130
rect 2475 -2506 2509 -130
rect 2653 -2506 2687 -130
rect 2831 -2506 2865 -130
rect 3009 -2506 3043 -130
rect 3187 -2506 3221 -130
rect 3365 -2506 3399 -130
rect 3543 -2506 3577 -130
rect 3721 -2506 3755 -130
rect 3899 -2506 3933 -130
rect 4077 -2506 4111 -130
rect 4255 -2506 4289 -130
rect 4433 -2506 4467 -130
rect 4611 -2506 4645 -130
rect 4789 -2506 4823 -130
rect 4967 -2506 5001 -130
rect 5145 -2506 5179 -130
rect 5323 -2506 5357 -130
rect 5501 -2506 5535 -130
rect 5679 -2506 5713 -130
rect 5857 -2506 5891 -130
rect 6035 -2506 6069 -130
rect 6213 -2506 6247 -130
rect 6391 -2506 6425 -130
rect 6569 -2506 6603 -130
rect 6747 -2506 6781 -130
rect 6925 -2506 6959 -130
rect 7103 -2506 7137 -130
rect 7281 -2506 7315 -130
rect 7459 -2506 7493 -130
rect 7637 -2506 7671 -130
rect 7815 -2506 7849 -130
rect 7993 -2506 8027 -130
rect 8171 -2506 8205 -130
rect 8349 -2506 8383 -130
rect 8527 -2506 8561 -130
rect 8705 -2506 8739 -130
rect 8883 -2506 8917 -130
<< nsubdiff >>
rect -9031 2667 -8935 2701
rect 8935 2667 9031 2701
rect -9031 2605 -8997 2667
rect 8997 2605 9031 2667
rect -9031 -2667 -8997 -2605
rect 8997 -2667 9031 -2605
rect -9031 -2701 -8935 -2667
rect 8935 -2701 9031 -2667
<< nsubdiffcont >>
rect -8935 2667 8935 2701
rect -9031 -2605 -8997 2605
rect 8997 -2605 9031 2605
rect -8935 -2701 8935 -2667
<< poly >>
rect -8871 2599 -8751 2615
rect -8871 2565 -8855 2599
rect -8767 2565 -8751 2599
rect -8871 2518 -8751 2565
rect -8693 2599 -8573 2615
rect -8693 2565 -8677 2599
rect -8589 2565 -8573 2599
rect -8693 2518 -8573 2565
rect -8515 2599 -8395 2615
rect -8515 2565 -8499 2599
rect -8411 2565 -8395 2599
rect -8515 2518 -8395 2565
rect -8337 2599 -8217 2615
rect -8337 2565 -8321 2599
rect -8233 2565 -8217 2599
rect -8337 2518 -8217 2565
rect -8159 2599 -8039 2615
rect -8159 2565 -8143 2599
rect -8055 2565 -8039 2599
rect -8159 2518 -8039 2565
rect -7981 2599 -7861 2615
rect -7981 2565 -7965 2599
rect -7877 2565 -7861 2599
rect -7981 2518 -7861 2565
rect -7803 2599 -7683 2615
rect -7803 2565 -7787 2599
rect -7699 2565 -7683 2599
rect -7803 2518 -7683 2565
rect -7625 2599 -7505 2615
rect -7625 2565 -7609 2599
rect -7521 2565 -7505 2599
rect -7625 2518 -7505 2565
rect -7447 2599 -7327 2615
rect -7447 2565 -7431 2599
rect -7343 2565 -7327 2599
rect -7447 2518 -7327 2565
rect -7269 2599 -7149 2615
rect -7269 2565 -7253 2599
rect -7165 2565 -7149 2599
rect -7269 2518 -7149 2565
rect -7091 2599 -6971 2615
rect -7091 2565 -7075 2599
rect -6987 2565 -6971 2599
rect -7091 2518 -6971 2565
rect -6913 2599 -6793 2615
rect -6913 2565 -6897 2599
rect -6809 2565 -6793 2599
rect -6913 2518 -6793 2565
rect -6735 2599 -6615 2615
rect -6735 2565 -6719 2599
rect -6631 2565 -6615 2599
rect -6735 2518 -6615 2565
rect -6557 2599 -6437 2615
rect -6557 2565 -6541 2599
rect -6453 2565 -6437 2599
rect -6557 2518 -6437 2565
rect -6379 2599 -6259 2615
rect -6379 2565 -6363 2599
rect -6275 2565 -6259 2599
rect -6379 2518 -6259 2565
rect -6201 2599 -6081 2615
rect -6201 2565 -6185 2599
rect -6097 2565 -6081 2599
rect -6201 2518 -6081 2565
rect -6023 2599 -5903 2615
rect -6023 2565 -6007 2599
rect -5919 2565 -5903 2599
rect -6023 2518 -5903 2565
rect -5845 2599 -5725 2615
rect -5845 2565 -5829 2599
rect -5741 2565 -5725 2599
rect -5845 2518 -5725 2565
rect -5667 2599 -5547 2615
rect -5667 2565 -5651 2599
rect -5563 2565 -5547 2599
rect -5667 2518 -5547 2565
rect -5489 2599 -5369 2615
rect -5489 2565 -5473 2599
rect -5385 2565 -5369 2599
rect -5489 2518 -5369 2565
rect -5311 2599 -5191 2615
rect -5311 2565 -5295 2599
rect -5207 2565 -5191 2599
rect -5311 2518 -5191 2565
rect -5133 2599 -5013 2615
rect -5133 2565 -5117 2599
rect -5029 2565 -5013 2599
rect -5133 2518 -5013 2565
rect -4955 2599 -4835 2615
rect -4955 2565 -4939 2599
rect -4851 2565 -4835 2599
rect -4955 2518 -4835 2565
rect -4777 2599 -4657 2615
rect -4777 2565 -4761 2599
rect -4673 2565 -4657 2599
rect -4777 2518 -4657 2565
rect -4599 2599 -4479 2615
rect -4599 2565 -4583 2599
rect -4495 2565 -4479 2599
rect -4599 2518 -4479 2565
rect -4421 2599 -4301 2615
rect -4421 2565 -4405 2599
rect -4317 2565 -4301 2599
rect -4421 2518 -4301 2565
rect -4243 2599 -4123 2615
rect -4243 2565 -4227 2599
rect -4139 2565 -4123 2599
rect -4243 2518 -4123 2565
rect -4065 2599 -3945 2615
rect -4065 2565 -4049 2599
rect -3961 2565 -3945 2599
rect -4065 2518 -3945 2565
rect -3887 2599 -3767 2615
rect -3887 2565 -3871 2599
rect -3783 2565 -3767 2599
rect -3887 2518 -3767 2565
rect -3709 2599 -3589 2615
rect -3709 2565 -3693 2599
rect -3605 2565 -3589 2599
rect -3709 2518 -3589 2565
rect -3531 2599 -3411 2615
rect -3531 2565 -3515 2599
rect -3427 2565 -3411 2599
rect -3531 2518 -3411 2565
rect -3353 2599 -3233 2615
rect -3353 2565 -3337 2599
rect -3249 2565 -3233 2599
rect -3353 2518 -3233 2565
rect -3175 2599 -3055 2615
rect -3175 2565 -3159 2599
rect -3071 2565 -3055 2599
rect -3175 2518 -3055 2565
rect -2997 2599 -2877 2615
rect -2997 2565 -2981 2599
rect -2893 2565 -2877 2599
rect -2997 2518 -2877 2565
rect -2819 2599 -2699 2615
rect -2819 2565 -2803 2599
rect -2715 2565 -2699 2599
rect -2819 2518 -2699 2565
rect -2641 2599 -2521 2615
rect -2641 2565 -2625 2599
rect -2537 2565 -2521 2599
rect -2641 2518 -2521 2565
rect -2463 2599 -2343 2615
rect -2463 2565 -2447 2599
rect -2359 2565 -2343 2599
rect -2463 2518 -2343 2565
rect -2285 2599 -2165 2615
rect -2285 2565 -2269 2599
rect -2181 2565 -2165 2599
rect -2285 2518 -2165 2565
rect -2107 2599 -1987 2615
rect -2107 2565 -2091 2599
rect -2003 2565 -1987 2599
rect -2107 2518 -1987 2565
rect -1929 2599 -1809 2615
rect -1929 2565 -1913 2599
rect -1825 2565 -1809 2599
rect -1929 2518 -1809 2565
rect -1751 2599 -1631 2615
rect -1751 2565 -1735 2599
rect -1647 2565 -1631 2599
rect -1751 2518 -1631 2565
rect -1573 2599 -1453 2615
rect -1573 2565 -1557 2599
rect -1469 2565 -1453 2599
rect -1573 2518 -1453 2565
rect -1395 2599 -1275 2615
rect -1395 2565 -1379 2599
rect -1291 2565 -1275 2599
rect -1395 2518 -1275 2565
rect -1217 2599 -1097 2615
rect -1217 2565 -1201 2599
rect -1113 2565 -1097 2599
rect -1217 2518 -1097 2565
rect -1039 2599 -919 2615
rect -1039 2565 -1023 2599
rect -935 2565 -919 2599
rect -1039 2518 -919 2565
rect -861 2599 -741 2615
rect -861 2565 -845 2599
rect -757 2565 -741 2599
rect -861 2518 -741 2565
rect -683 2599 -563 2615
rect -683 2565 -667 2599
rect -579 2565 -563 2599
rect -683 2518 -563 2565
rect -505 2599 -385 2615
rect -505 2565 -489 2599
rect -401 2565 -385 2599
rect -505 2518 -385 2565
rect -327 2599 -207 2615
rect -327 2565 -311 2599
rect -223 2565 -207 2599
rect -327 2518 -207 2565
rect -149 2599 -29 2615
rect -149 2565 -133 2599
rect -45 2565 -29 2599
rect -149 2518 -29 2565
rect 29 2599 149 2615
rect 29 2565 45 2599
rect 133 2565 149 2599
rect 29 2518 149 2565
rect 207 2599 327 2615
rect 207 2565 223 2599
rect 311 2565 327 2599
rect 207 2518 327 2565
rect 385 2599 505 2615
rect 385 2565 401 2599
rect 489 2565 505 2599
rect 385 2518 505 2565
rect 563 2599 683 2615
rect 563 2565 579 2599
rect 667 2565 683 2599
rect 563 2518 683 2565
rect 741 2599 861 2615
rect 741 2565 757 2599
rect 845 2565 861 2599
rect 741 2518 861 2565
rect 919 2599 1039 2615
rect 919 2565 935 2599
rect 1023 2565 1039 2599
rect 919 2518 1039 2565
rect 1097 2599 1217 2615
rect 1097 2565 1113 2599
rect 1201 2565 1217 2599
rect 1097 2518 1217 2565
rect 1275 2599 1395 2615
rect 1275 2565 1291 2599
rect 1379 2565 1395 2599
rect 1275 2518 1395 2565
rect 1453 2599 1573 2615
rect 1453 2565 1469 2599
rect 1557 2565 1573 2599
rect 1453 2518 1573 2565
rect 1631 2599 1751 2615
rect 1631 2565 1647 2599
rect 1735 2565 1751 2599
rect 1631 2518 1751 2565
rect 1809 2599 1929 2615
rect 1809 2565 1825 2599
rect 1913 2565 1929 2599
rect 1809 2518 1929 2565
rect 1987 2599 2107 2615
rect 1987 2565 2003 2599
rect 2091 2565 2107 2599
rect 1987 2518 2107 2565
rect 2165 2599 2285 2615
rect 2165 2565 2181 2599
rect 2269 2565 2285 2599
rect 2165 2518 2285 2565
rect 2343 2599 2463 2615
rect 2343 2565 2359 2599
rect 2447 2565 2463 2599
rect 2343 2518 2463 2565
rect 2521 2599 2641 2615
rect 2521 2565 2537 2599
rect 2625 2565 2641 2599
rect 2521 2518 2641 2565
rect 2699 2599 2819 2615
rect 2699 2565 2715 2599
rect 2803 2565 2819 2599
rect 2699 2518 2819 2565
rect 2877 2599 2997 2615
rect 2877 2565 2893 2599
rect 2981 2565 2997 2599
rect 2877 2518 2997 2565
rect 3055 2599 3175 2615
rect 3055 2565 3071 2599
rect 3159 2565 3175 2599
rect 3055 2518 3175 2565
rect 3233 2599 3353 2615
rect 3233 2565 3249 2599
rect 3337 2565 3353 2599
rect 3233 2518 3353 2565
rect 3411 2599 3531 2615
rect 3411 2565 3427 2599
rect 3515 2565 3531 2599
rect 3411 2518 3531 2565
rect 3589 2599 3709 2615
rect 3589 2565 3605 2599
rect 3693 2565 3709 2599
rect 3589 2518 3709 2565
rect 3767 2599 3887 2615
rect 3767 2565 3783 2599
rect 3871 2565 3887 2599
rect 3767 2518 3887 2565
rect 3945 2599 4065 2615
rect 3945 2565 3961 2599
rect 4049 2565 4065 2599
rect 3945 2518 4065 2565
rect 4123 2599 4243 2615
rect 4123 2565 4139 2599
rect 4227 2565 4243 2599
rect 4123 2518 4243 2565
rect 4301 2599 4421 2615
rect 4301 2565 4317 2599
rect 4405 2565 4421 2599
rect 4301 2518 4421 2565
rect 4479 2599 4599 2615
rect 4479 2565 4495 2599
rect 4583 2565 4599 2599
rect 4479 2518 4599 2565
rect 4657 2599 4777 2615
rect 4657 2565 4673 2599
rect 4761 2565 4777 2599
rect 4657 2518 4777 2565
rect 4835 2599 4955 2615
rect 4835 2565 4851 2599
rect 4939 2565 4955 2599
rect 4835 2518 4955 2565
rect 5013 2599 5133 2615
rect 5013 2565 5029 2599
rect 5117 2565 5133 2599
rect 5013 2518 5133 2565
rect 5191 2599 5311 2615
rect 5191 2565 5207 2599
rect 5295 2565 5311 2599
rect 5191 2518 5311 2565
rect 5369 2599 5489 2615
rect 5369 2565 5385 2599
rect 5473 2565 5489 2599
rect 5369 2518 5489 2565
rect 5547 2599 5667 2615
rect 5547 2565 5563 2599
rect 5651 2565 5667 2599
rect 5547 2518 5667 2565
rect 5725 2599 5845 2615
rect 5725 2565 5741 2599
rect 5829 2565 5845 2599
rect 5725 2518 5845 2565
rect 5903 2599 6023 2615
rect 5903 2565 5919 2599
rect 6007 2565 6023 2599
rect 5903 2518 6023 2565
rect 6081 2599 6201 2615
rect 6081 2565 6097 2599
rect 6185 2565 6201 2599
rect 6081 2518 6201 2565
rect 6259 2599 6379 2615
rect 6259 2565 6275 2599
rect 6363 2565 6379 2599
rect 6259 2518 6379 2565
rect 6437 2599 6557 2615
rect 6437 2565 6453 2599
rect 6541 2565 6557 2599
rect 6437 2518 6557 2565
rect 6615 2599 6735 2615
rect 6615 2565 6631 2599
rect 6719 2565 6735 2599
rect 6615 2518 6735 2565
rect 6793 2599 6913 2615
rect 6793 2565 6809 2599
rect 6897 2565 6913 2599
rect 6793 2518 6913 2565
rect 6971 2599 7091 2615
rect 6971 2565 6987 2599
rect 7075 2565 7091 2599
rect 6971 2518 7091 2565
rect 7149 2599 7269 2615
rect 7149 2565 7165 2599
rect 7253 2565 7269 2599
rect 7149 2518 7269 2565
rect 7327 2599 7447 2615
rect 7327 2565 7343 2599
rect 7431 2565 7447 2599
rect 7327 2518 7447 2565
rect 7505 2599 7625 2615
rect 7505 2565 7521 2599
rect 7609 2565 7625 2599
rect 7505 2518 7625 2565
rect 7683 2599 7803 2615
rect 7683 2565 7699 2599
rect 7787 2565 7803 2599
rect 7683 2518 7803 2565
rect 7861 2599 7981 2615
rect 7861 2565 7877 2599
rect 7965 2565 7981 2599
rect 7861 2518 7981 2565
rect 8039 2599 8159 2615
rect 8039 2565 8055 2599
rect 8143 2565 8159 2599
rect 8039 2518 8159 2565
rect 8217 2599 8337 2615
rect 8217 2565 8233 2599
rect 8321 2565 8337 2599
rect 8217 2518 8337 2565
rect 8395 2599 8515 2615
rect 8395 2565 8411 2599
rect 8499 2565 8515 2599
rect 8395 2518 8515 2565
rect 8573 2599 8693 2615
rect 8573 2565 8589 2599
rect 8677 2565 8693 2599
rect 8573 2518 8693 2565
rect 8751 2599 8871 2615
rect 8751 2565 8767 2599
rect 8855 2565 8871 2599
rect 8751 2518 8871 2565
rect -8871 71 -8751 118
rect -8871 37 -8855 71
rect -8767 37 -8751 71
rect -8871 21 -8751 37
rect -8693 71 -8573 118
rect -8693 37 -8677 71
rect -8589 37 -8573 71
rect -8693 21 -8573 37
rect -8515 71 -8395 118
rect -8515 37 -8499 71
rect -8411 37 -8395 71
rect -8515 21 -8395 37
rect -8337 71 -8217 118
rect -8337 37 -8321 71
rect -8233 37 -8217 71
rect -8337 21 -8217 37
rect -8159 71 -8039 118
rect -8159 37 -8143 71
rect -8055 37 -8039 71
rect -8159 21 -8039 37
rect -7981 71 -7861 118
rect -7981 37 -7965 71
rect -7877 37 -7861 71
rect -7981 21 -7861 37
rect -7803 71 -7683 118
rect -7803 37 -7787 71
rect -7699 37 -7683 71
rect -7803 21 -7683 37
rect -7625 71 -7505 118
rect -7625 37 -7609 71
rect -7521 37 -7505 71
rect -7625 21 -7505 37
rect -7447 71 -7327 118
rect -7447 37 -7431 71
rect -7343 37 -7327 71
rect -7447 21 -7327 37
rect -7269 71 -7149 118
rect -7269 37 -7253 71
rect -7165 37 -7149 71
rect -7269 21 -7149 37
rect -7091 71 -6971 118
rect -7091 37 -7075 71
rect -6987 37 -6971 71
rect -7091 21 -6971 37
rect -6913 71 -6793 118
rect -6913 37 -6897 71
rect -6809 37 -6793 71
rect -6913 21 -6793 37
rect -6735 71 -6615 118
rect -6735 37 -6719 71
rect -6631 37 -6615 71
rect -6735 21 -6615 37
rect -6557 71 -6437 118
rect -6557 37 -6541 71
rect -6453 37 -6437 71
rect -6557 21 -6437 37
rect -6379 71 -6259 118
rect -6379 37 -6363 71
rect -6275 37 -6259 71
rect -6379 21 -6259 37
rect -6201 71 -6081 118
rect -6201 37 -6185 71
rect -6097 37 -6081 71
rect -6201 21 -6081 37
rect -6023 71 -5903 118
rect -6023 37 -6007 71
rect -5919 37 -5903 71
rect -6023 21 -5903 37
rect -5845 71 -5725 118
rect -5845 37 -5829 71
rect -5741 37 -5725 71
rect -5845 21 -5725 37
rect -5667 71 -5547 118
rect -5667 37 -5651 71
rect -5563 37 -5547 71
rect -5667 21 -5547 37
rect -5489 71 -5369 118
rect -5489 37 -5473 71
rect -5385 37 -5369 71
rect -5489 21 -5369 37
rect -5311 71 -5191 118
rect -5311 37 -5295 71
rect -5207 37 -5191 71
rect -5311 21 -5191 37
rect -5133 71 -5013 118
rect -5133 37 -5117 71
rect -5029 37 -5013 71
rect -5133 21 -5013 37
rect -4955 71 -4835 118
rect -4955 37 -4939 71
rect -4851 37 -4835 71
rect -4955 21 -4835 37
rect -4777 71 -4657 118
rect -4777 37 -4761 71
rect -4673 37 -4657 71
rect -4777 21 -4657 37
rect -4599 71 -4479 118
rect -4599 37 -4583 71
rect -4495 37 -4479 71
rect -4599 21 -4479 37
rect -4421 71 -4301 118
rect -4421 37 -4405 71
rect -4317 37 -4301 71
rect -4421 21 -4301 37
rect -4243 71 -4123 118
rect -4243 37 -4227 71
rect -4139 37 -4123 71
rect -4243 21 -4123 37
rect -4065 71 -3945 118
rect -4065 37 -4049 71
rect -3961 37 -3945 71
rect -4065 21 -3945 37
rect -3887 71 -3767 118
rect -3887 37 -3871 71
rect -3783 37 -3767 71
rect -3887 21 -3767 37
rect -3709 71 -3589 118
rect -3709 37 -3693 71
rect -3605 37 -3589 71
rect -3709 21 -3589 37
rect -3531 71 -3411 118
rect -3531 37 -3515 71
rect -3427 37 -3411 71
rect -3531 21 -3411 37
rect -3353 71 -3233 118
rect -3353 37 -3337 71
rect -3249 37 -3233 71
rect -3353 21 -3233 37
rect -3175 71 -3055 118
rect -3175 37 -3159 71
rect -3071 37 -3055 71
rect -3175 21 -3055 37
rect -2997 71 -2877 118
rect -2997 37 -2981 71
rect -2893 37 -2877 71
rect -2997 21 -2877 37
rect -2819 71 -2699 118
rect -2819 37 -2803 71
rect -2715 37 -2699 71
rect -2819 21 -2699 37
rect -2641 71 -2521 118
rect -2641 37 -2625 71
rect -2537 37 -2521 71
rect -2641 21 -2521 37
rect -2463 71 -2343 118
rect -2463 37 -2447 71
rect -2359 37 -2343 71
rect -2463 21 -2343 37
rect -2285 71 -2165 118
rect -2285 37 -2269 71
rect -2181 37 -2165 71
rect -2285 21 -2165 37
rect -2107 71 -1987 118
rect -2107 37 -2091 71
rect -2003 37 -1987 71
rect -2107 21 -1987 37
rect -1929 71 -1809 118
rect -1929 37 -1913 71
rect -1825 37 -1809 71
rect -1929 21 -1809 37
rect -1751 71 -1631 118
rect -1751 37 -1735 71
rect -1647 37 -1631 71
rect -1751 21 -1631 37
rect -1573 71 -1453 118
rect -1573 37 -1557 71
rect -1469 37 -1453 71
rect -1573 21 -1453 37
rect -1395 71 -1275 118
rect -1395 37 -1379 71
rect -1291 37 -1275 71
rect -1395 21 -1275 37
rect -1217 71 -1097 118
rect -1217 37 -1201 71
rect -1113 37 -1097 71
rect -1217 21 -1097 37
rect -1039 71 -919 118
rect -1039 37 -1023 71
rect -935 37 -919 71
rect -1039 21 -919 37
rect -861 71 -741 118
rect -861 37 -845 71
rect -757 37 -741 71
rect -861 21 -741 37
rect -683 71 -563 118
rect -683 37 -667 71
rect -579 37 -563 71
rect -683 21 -563 37
rect -505 71 -385 118
rect -505 37 -489 71
rect -401 37 -385 71
rect -505 21 -385 37
rect -327 71 -207 118
rect -327 37 -311 71
rect -223 37 -207 71
rect -327 21 -207 37
rect -149 71 -29 118
rect -149 37 -133 71
rect -45 37 -29 71
rect -149 21 -29 37
rect 29 71 149 118
rect 29 37 45 71
rect 133 37 149 71
rect 29 21 149 37
rect 207 71 327 118
rect 207 37 223 71
rect 311 37 327 71
rect 207 21 327 37
rect 385 71 505 118
rect 385 37 401 71
rect 489 37 505 71
rect 385 21 505 37
rect 563 71 683 118
rect 563 37 579 71
rect 667 37 683 71
rect 563 21 683 37
rect 741 71 861 118
rect 741 37 757 71
rect 845 37 861 71
rect 741 21 861 37
rect 919 71 1039 118
rect 919 37 935 71
rect 1023 37 1039 71
rect 919 21 1039 37
rect 1097 71 1217 118
rect 1097 37 1113 71
rect 1201 37 1217 71
rect 1097 21 1217 37
rect 1275 71 1395 118
rect 1275 37 1291 71
rect 1379 37 1395 71
rect 1275 21 1395 37
rect 1453 71 1573 118
rect 1453 37 1469 71
rect 1557 37 1573 71
rect 1453 21 1573 37
rect 1631 71 1751 118
rect 1631 37 1647 71
rect 1735 37 1751 71
rect 1631 21 1751 37
rect 1809 71 1929 118
rect 1809 37 1825 71
rect 1913 37 1929 71
rect 1809 21 1929 37
rect 1987 71 2107 118
rect 1987 37 2003 71
rect 2091 37 2107 71
rect 1987 21 2107 37
rect 2165 71 2285 118
rect 2165 37 2181 71
rect 2269 37 2285 71
rect 2165 21 2285 37
rect 2343 71 2463 118
rect 2343 37 2359 71
rect 2447 37 2463 71
rect 2343 21 2463 37
rect 2521 71 2641 118
rect 2521 37 2537 71
rect 2625 37 2641 71
rect 2521 21 2641 37
rect 2699 71 2819 118
rect 2699 37 2715 71
rect 2803 37 2819 71
rect 2699 21 2819 37
rect 2877 71 2997 118
rect 2877 37 2893 71
rect 2981 37 2997 71
rect 2877 21 2997 37
rect 3055 71 3175 118
rect 3055 37 3071 71
rect 3159 37 3175 71
rect 3055 21 3175 37
rect 3233 71 3353 118
rect 3233 37 3249 71
rect 3337 37 3353 71
rect 3233 21 3353 37
rect 3411 71 3531 118
rect 3411 37 3427 71
rect 3515 37 3531 71
rect 3411 21 3531 37
rect 3589 71 3709 118
rect 3589 37 3605 71
rect 3693 37 3709 71
rect 3589 21 3709 37
rect 3767 71 3887 118
rect 3767 37 3783 71
rect 3871 37 3887 71
rect 3767 21 3887 37
rect 3945 71 4065 118
rect 3945 37 3961 71
rect 4049 37 4065 71
rect 3945 21 4065 37
rect 4123 71 4243 118
rect 4123 37 4139 71
rect 4227 37 4243 71
rect 4123 21 4243 37
rect 4301 71 4421 118
rect 4301 37 4317 71
rect 4405 37 4421 71
rect 4301 21 4421 37
rect 4479 71 4599 118
rect 4479 37 4495 71
rect 4583 37 4599 71
rect 4479 21 4599 37
rect 4657 71 4777 118
rect 4657 37 4673 71
rect 4761 37 4777 71
rect 4657 21 4777 37
rect 4835 71 4955 118
rect 4835 37 4851 71
rect 4939 37 4955 71
rect 4835 21 4955 37
rect 5013 71 5133 118
rect 5013 37 5029 71
rect 5117 37 5133 71
rect 5013 21 5133 37
rect 5191 71 5311 118
rect 5191 37 5207 71
rect 5295 37 5311 71
rect 5191 21 5311 37
rect 5369 71 5489 118
rect 5369 37 5385 71
rect 5473 37 5489 71
rect 5369 21 5489 37
rect 5547 71 5667 118
rect 5547 37 5563 71
rect 5651 37 5667 71
rect 5547 21 5667 37
rect 5725 71 5845 118
rect 5725 37 5741 71
rect 5829 37 5845 71
rect 5725 21 5845 37
rect 5903 71 6023 118
rect 5903 37 5919 71
rect 6007 37 6023 71
rect 5903 21 6023 37
rect 6081 71 6201 118
rect 6081 37 6097 71
rect 6185 37 6201 71
rect 6081 21 6201 37
rect 6259 71 6379 118
rect 6259 37 6275 71
rect 6363 37 6379 71
rect 6259 21 6379 37
rect 6437 71 6557 118
rect 6437 37 6453 71
rect 6541 37 6557 71
rect 6437 21 6557 37
rect 6615 71 6735 118
rect 6615 37 6631 71
rect 6719 37 6735 71
rect 6615 21 6735 37
rect 6793 71 6913 118
rect 6793 37 6809 71
rect 6897 37 6913 71
rect 6793 21 6913 37
rect 6971 71 7091 118
rect 6971 37 6987 71
rect 7075 37 7091 71
rect 6971 21 7091 37
rect 7149 71 7269 118
rect 7149 37 7165 71
rect 7253 37 7269 71
rect 7149 21 7269 37
rect 7327 71 7447 118
rect 7327 37 7343 71
rect 7431 37 7447 71
rect 7327 21 7447 37
rect 7505 71 7625 118
rect 7505 37 7521 71
rect 7609 37 7625 71
rect 7505 21 7625 37
rect 7683 71 7803 118
rect 7683 37 7699 71
rect 7787 37 7803 71
rect 7683 21 7803 37
rect 7861 71 7981 118
rect 7861 37 7877 71
rect 7965 37 7981 71
rect 7861 21 7981 37
rect 8039 71 8159 118
rect 8039 37 8055 71
rect 8143 37 8159 71
rect 8039 21 8159 37
rect 8217 71 8337 118
rect 8217 37 8233 71
rect 8321 37 8337 71
rect 8217 21 8337 37
rect 8395 71 8515 118
rect 8395 37 8411 71
rect 8499 37 8515 71
rect 8395 21 8515 37
rect 8573 71 8693 118
rect 8573 37 8589 71
rect 8677 37 8693 71
rect 8573 21 8693 37
rect 8751 71 8871 118
rect 8751 37 8767 71
rect 8855 37 8871 71
rect 8751 21 8871 37
rect -8871 -37 -8751 -21
rect -8871 -71 -8855 -37
rect -8767 -71 -8751 -37
rect -8871 -118 -8751 -71
rect -8693 -37 -8573 -21
rect -8693 -71 -8677 -37
rect -8589 -71 -8573 -37
rect -8693 -118 -8573 -71
rect -8515 -37 -8395 -21
rect -8515 -71 -8499 -37
rect -8411 -71 -8395 -37
rect -8515 -118 -8395 -71
rect -8337 -37 -8217 -21
rect -8337 -71 -8321 -37
rect -8233 -71 -8217 -37
rect -8337 -118 -8217 -71
rect -8159 -37 -8039 -21
rect -8159 -71 -8143 -37
rect -8055 -71 -8039 -37
rect -8159 -118 -8039 -71
rect -7981 -37 -7861 -21
rect -7981 -71 -7965 -37
rect -7877 -71 -7861 -37
rect -7981 -118 -7861 -71
rect -7803 -37 -7683 -21
rect -7803 -71 -7787 -37
rect -7699 -71 -7683 -37
rect -7803 -118 -7683 -71
rect -7625 -37 -7505 -21
rect -7625 -71 -7609 -37
rect -7521 -71 -7505 -37
rect -7625 -118 -7505 -71
rect -7447 -37 -7327 -21
rect -7447 -71 -7431 -37
rect -7343 -71 -7327 -37
rect -7447 -118 -7327 -71
rect -7269 -37 -7149 -21
rect -7269 -71 -7253 -37
rect -7165 -71 -7149 -37
rect -7269 -118 -7149 -71
rect -7091 -37 -6971 -21
rect -7091 -71 -7075 -37
rect -6987 -71 -6971 -37
rect -7091 -118 -6971 -71
rect -6913 -37 -6793 -21
rect -6913 -71 -6897 -37
rect -6809 -71 -6793 -37
rect -6913 -118 -6793 -71
rect -6735 -37 -6615 -21
rect -6735 -71 -6719 -37
rect -6631 -71 -6615 -37
rect -6735 -118 -6615 -71
rect -6557 -37 -6437 -21
rect -6557 -71 -6541 -37
rect -6453 -71 -6437 -37
rect -6557 -118 -6437 -71
rect -6379 -37 -6259 -21
rect -6379 -71 -6363 -37
rect -6275 -71 -6259 -37
rect -6379 -118 -6259 -71
rect -6201 -37 -6081 -21
rect -6201 -71 -6185 -37
rect -6097 -71 -6081 -37
rect -6201 -118 -6081 -71
rect -6023 -37 -5903 -21
rect -6023 -71 -6007 -37
rect -5919 -71 -5903 -37
rect -6023 -118 -5903 -71
rect -5845 -37 -5725 -21
rect -5845 -71 -5829 -37
rect -5741 -71 -5725 -37
rect -5845 -118 -5725 -71
rect -5667 -37 -5547 -21
rect -5667 -71 -5651 -37
rect -5563 -71 -5547 -37
rect -5667 -118 -5547 -71
rect -5489 -37 -5369 -21
rect -5489 -71 -5473 -37
rect -5385 -71 -5369 -37
rect -5489 -118 -5369 -71
rect -5311 -37 -5191 -21
rect -5311 -71 -5295 -37
rect -5207 -71 -5191 -37
rect -5311 -118 -5191 -71
rect -5133 -37 -5013 -21
rect -5133 -71 -5117 -37
rect -5029 -71 -5013 -37
rect -5133 -118 -5013 -71
rect -4955 -37 -4835 -21
rect -4955 -71 -4939 -37
rect -4851 -71 -4835 -37
rect -4955 -118 -4835 -71
rect -4777 -37 -4657 -21
rect -4777 -71 -4761 -37
rect -4673 -71 -4657 -37
rect -4777 -118 -4657 -71
rect -4599 -37 -4479 -21
rect -4599 -71 -4583 -37
rect -4495 -71 -4479 -37
rect -4599 -118 -4479 -71
rect -4421 -37 -4301 -21
rect -4421 -71 -4405 -37
rect -4317 -71 -4301 -37
rect -4421 -118 -4301 -71
rect -4243 -37 -4123 -21
rect -4243 -71 -4227 -37
rect -4139 -71 -4123 -37
rect -4243 -118 -4123 -71
rect -4065 -37 -3945 -21
rect -4065 -71 -4049 -37
rect -3961 -71 -3945 -37
rect -4065 -118 -3945 -71
rect -3887 -37 -3767 -21
rect -3887 -71 -3871 -37
rect -3783 -71 -3767 -37
rect -3887 -118 -3767 -71
rect -3709 -37 -3589 -21
rect -3709 -71 -3693 -37
rect -3605 -71 -3589 -37
rect -3709 -118 -3589 -71
rect -3531 -37 -3411 -21
rect -3531 -71 -3515 -37
rect -3427 -71 -3411 -37
rect -3531 -118 -3411 -71
rect -3353 -37 -3233 -21
rect -3353 -71 -3337 -37
rect -3249 -71 -3233 -37
rect -3353 -118 -3233 -71
rect -3175 -37 -3055 -21
rect -3175 -71 -3159 -37
rect -3071 -71 -3055 -37
rect -3175 -118 -3055 -71
rect -2997 -37 -2877 -21
rect -2997 -71 -2981 -37
rect -2893 -71 -2877 -37
rect -2997 -118 -2877 -71
rect -2819 -37 -2699 -21
rect -2819 -71 -2803 -37
rect -2715 -71 -2699 -37
rect -2819 -118 -2699 -71
rect -2641 -37 -2521 -21
rect -2641 -71 -2625 -37
rect -2537 -71 -2521 -37
rect -2641 -118 -2521 -71
rect -2463 -37 -2343 -21
rect -2463 -71 -2447 -37
rect -2359 -71 -2343 -37
rect -2463 -118 -2343 -71
rect -2285 -37 -2165 -21
rect -2285 -71 -2269 -37
rect -2181 -71 -2165 -37
rect -2285 -118 -2165 -71
rect -2107 -37 -1987 -21
rect -2107 -71 -2091 -37
rect -2003 -71 -1987 -37
rect -2107 -118 -1987 -71
rect -1929 -37 -1809 -21
rect -1929 -71 -1913 -37
rect -1825 -71 -1809 -37
rect -1929 -118 -1809 -71
rect -1751 -37 -1631 -21
rect -1751 -71 -1735 -37
rect -1647 -71 -1631 -37
rect -1751 -118 -1631 -71
rect -1573 -37 -1453 -21
rect -1573 -71 -1557 -37
rect -1469 -71 -1453 -37
rect -1573 -118 -1453 -71
rect -1395 -37 -1275 -21
rect -1395 -71 -1379 -37
rect -1291 -71 -1275 -37
rect -1395 -118 -1275 -71
rect -1217 -37 -1097 -21
rect -1217 -71 -1201 -37
rect -1113 -71 -1097 -37
rect -1217 -118 -1097 -71
rect -1039 -37 -919 -21
rect -1039 -71 -1023 -37
rect -935 -71 -919 -37
rect -1039 -118 -919 -71
rect -861 -37 -741 -21
rect -861 -71 -845 -37
rect -757 -71 -741 -37
rect -861 -118 -741 -71
rect -683 -37 -563 -21
rect -683 -71 -667 -37
rect -579 -71 -563 -37
rect -683 -118 -563 -71
rect -505 -37 -385 -21
rect -505 -71 -489 -37
rect -401 -71 -385 -37
rect -505 -118 -385 -71
rect -327 -37 -207 -21
rect -327 -71 -311 -37
rect -223 -71 -207 -37
rect -327 -118 -207 -71
rect -149 -37 -29 -21
rect -149 -71 -133 -37
rect -45 -71 -29 -37
rect -149 -118 -29 -71
rect 29 -37 149 -21
rect 29 -71 45 -37
rect 133 -71 149 -37
rect 29 -118 149 -71
rect 207 -37 327 -21
rect 207 -71 223 -37
rect 311 -71 327 -37
rect 207 -118 327 -71
rect 385 -37 505 -21
rect 385 -71 401 -37
rect 489 -71 505 -37
rect 385 -118 505 -71
rect 563 -37 683 -21
rect 563 -71 579 -37
rect 667 -71 683 -37
rect 563 -118 683 -71
rect 741 -37 861 -21
rect 741 -71 757 -37
rect 845 -71 861 -37
rect 741 -118 861 -71
rect 919 -37 1039 -21
rect 919 -71 935 -37
rect 1023 -71 1039 -37
rect 919 -118 1039 -71
rect 1097 -37 1217 -21
rect 1097 -71 1113 -37
rect 1201 -71 1217 -37
rect 1097 -118 1217 -71
rect 1275 -37 1395 -21
rect 1275 -71 1291 -37
rect 1379 -71 1395 -37
rect 1275 -118 1395 -71
rect 1453 -37 1573 -21
rect 1453 -71 1469 -37
rect 1557 -71 1573 -37
rect 1453 -118 1573 -71
rect 1631 -37 1751 -21
rect 1631 -71 1647 -37
rect 1735 -71 1751 -37
rect 1631 -118 1751 -71
rect 1809 -37 1929 -21
rect 1809 -71 1825 -37
rect 1913 -71 1929 -37
rect 1809 -118 1929 -71
rect 1987 -37 2107 -21
rect 1987 -71 2003 -37
rect 2091 -71 2107 -37
rect 1987 -118 2107 -71
rect 2165 -37 2285 -21
rect 2165 -71 2181 -37
rect 2269 -71 2285 -37
rect 2165 -118 2285 -71
rect 2343 -37 2463 -21
rect 2343 -71 2359 -37
rect 2447 -71 2463 -37
rect 2343 -118 2463 -71
rect 2521 -37 2641 -21
rect 2521 -71 2537 -37
rect 2625 -71 2641 -37
rect 2521 -118 2641 -71
rect 2699 -37 2819 -21
rect 2699 -71 2715 -37
rect 2803 -71 2819 -37
rect 2699 -118 2819 -71
rect 2877 -37 2997 -21
rect 2877 -71 2893 -37
rect 2981 -71 2997 -37
rect 2877 -118 2997 -71
rect 3055 -37 3175 -21
rect 3055 -71 3071 -37
rect 3159 -71 3175 -37
rect 3055 -118 3175 -71
rect 3233 -37 3353 -21
rect 3233 -71 3249 -37
rect 3337 -71 3353 -37
rect 3233 -118 3353 -71
rect 3411 -37 3531 -21
rect 3411 -71 3427 -37
rect 3515 -71 3531 -37
rect 3411 -118 3531 -71
rect 3589 -37 3709 -21
rect 3589 -71 3605 -37
rect 3693 -71 3709 -37
rect 3589 -118 3709 -71
rect 3767 -37 3887 -21
rect 3767 -71 3783 -37
rect 3871 -71 3887 -37
rect 3767 -118 3887 -71
rect 3945 -37 4065 -21
rect 3945 -71 3961 -37
rect 4049 -71 4065 -37
rect 3945 -118 4065 -71
rect 4123 -37 4243 -21
rect 4123 -71 4139 -37
rect 4227 -71 4243 -37
rect 4123 -118 4243 -71
rect 4301 -37 4421 -21
rect 4301 -71 4317 -37
rect 4405 -71 4421 -37
rect 4301 -118 4421 -71
rect 4479 -37 4599 -21
rect 4479 -71 4495 -37
rect 4583 -71 4599 -37
rect 4479 -118 4599 -71
rect 4657 -37 4777 -21
rect 4657 -71 4673 -37
rect 4761 -71 4777 -37
rect 4657 -118 4777 -71
rect 4835 -37 4955 -21
rect 4835 -71 4851 -37
rect 4939 -71 4955 -37
rect 4835 -118 4955 -71
rect 5013 -37 5133 -21
rect 5013 -71 5029 -37
rect 5117 -71 5133 -37
rect 5013 -118 5133 -71
rect 5191 -37 5311 -21
rect 5191 -71 5207 -37
rect 5295 -71 5311 -37
rect 5191 -118 5311 -71
rect 5369 -37 5489 -21
rect 5369 -71 5385 -37
rect 5473 -71 5489 -37
rect 5369 -118 5489 -71
rect 5547 -37 5667 -21
rect 5547 -71 5563 -37
rect 5651 -71 5667 -37
rect 5547 -118 5667 -71
rect 5725 -37 5845 -21
rect 5725 -71 5741 -37
rect 5829 -71 5845 -37
rect 5725 -118 5845 -71
rect 5903 -37 6023 -21
rect 5903 -71 5919 -37
rect 6007 -71 6023 -37
rect 5903 -118 6023 -71
rect 6081 -37 6201 -21
rect 6081 -71 6097 -37
rect 6185 -71 6201 -37
rect 6081 -118 6201 -71
rect 6259 -37 6379 -21
rect 6259 -71 6275 -37
rect 6363 -71 6379 -37
rect 6259 -118 6379 -71
rect 6437 -37 6557 -21
rect 6437 -71 6453 -37
rect 6541 -71 6557 -37
rect 6437 -118 6557 -71
rect 6615 -37 6735 -21
rect 6615 -71 6631 -37
rect 6719 -71 6735 -37
rect 6615 -118 6735 -71
rect 6793 -37 6913 -21
rect 6793 -71 6809 -37
rect 6897 -71 6913 -37
rect 6793 -118 6913 -71
rect 6971 -37 7091 -21
rect 6971 -71 6987 -37
rect 7075 -71 7091 -37
rect 6971 -118 7091 -71
rect 7149 -37 7269 -21
rect 7149 -71 7165 -37
rect 7253 -71 7269 -37
rect 7149 -118 7269 -71
rect 7327 -37 7447 -21
rect 7327 -71 7343 -37
rect 7431 -71 7447 -37
rect 7327 -118 7447 -71
rect 7505 -37 7625 -21
rect 7505 -71 7521 -37
rect 7609 -71 7625 -37
rect 7505 -118 7625 -71
rect 7683 -37 7803 -21
rect 7683 -71 7699 -37
rect 7787 -71 7803 -37
rect 7683 -118 7803 -71
rect 7861 -37 7981 -21
rect 7861 -71 7877 -37
rect 7965 -71 7981 -37
rect 7861 -118 7981 -71
rect 8039 -37 8159 -21
rect 8039 -71 8055 -37
rect 8143 -71 8159 -37
rect 8039 -118 8159 -71
rect 8217 -37 8337 -21
rect 8217 -71 8233 -37
rect 8321 -71 8337 -37
rect 8217 -118 8337 -71
rect 8395 -37 8515 -21
rect 8395 -71 8411 -37
rect 8499 -71 8515 -37
rect 8395 -118 8515 -71
rect 8573 -37 8693 -21
rect 8573 -71 8589 -37
rect 8677 -71 8693 -37
rect 8573 -118 8693 -71
rect 8751 -37 8871 -21
rect 8751 -71 8767 -37
rect 8855 -71 8871 -37
rect 8751 -118 8871 -71
rect -8871 -2565 -8751 -2518
rect -8871 -2599 -8855 -2565
rect -8767 -2599 -8751 -2565
rect -8871 -2615 -8751 -2599
rect -8693 -2565 -8573 -2518
rect -8693 -2599 -8677 -2565
rect -8589 -2599 -8573 -2565
rect -8693 -2615 -8573 -2599
rect -8515 -2565 -8395 -2518
rect -8515 -2599 -8499 -2565
rect -8411 -2599 -8395 -2565
rect -8515 -2615 -8395 -2599
rect -8337 -2565 -8217 -2518
rect -8337 -2599 -8321 -2565
rect -8233 -2599 -8217 -2565
rect -8337 -2615 -8217 -2599
rect -8159 -2565 -8039 -2518
rect -8159 -2599 -8143 -2565
rect -8055 -2599 -8039 -2565
rect -8159 -2615 -8039 -2599
rect -7981 -2565 -7861 -2518
rect -7981 -2599 -7965 -2565
rect -7877 -2599 -7861 -2565
rect -7981 -2615 -7861 -2599
rect -7803 -2565 -7683 -2518
rect -7803 -2599 -7787 -2565
rect -7699 -2599 -7683 -2565
rect -7803 -2615 -7683 -2599
rect -7625 -2565 -7505 -2518
rect -7625 -2599 -7609 -2565
rect -7521 -2599 -7505 -2565
rect -7625 -2615 -7505 -2599
rect -7447 -2565 -7327 -2518
rect -7447 -2599 -7431 -2565
rect -7343 -2599 -7327 -2565
rect -7447 -2615 -7327 -2599
rect -7269 -2565 -7149 -2518
rect -7269 -2599 -7253 -2565
rect -7165 -2599 -7149 -2565
rect -7269 -2615 -7149 -2599
rect -7091 -2565 -6971 -2518
rect -7091 -2599 -7075 -2565
rect -6987 -2599 -6971 -2565
rect -7091 -2615 -6971 -2599
rect -6913 -2565 -6793 -2518
rect -6913 -2599 -6897 -2565
rect -6809 -2599 -6793 -2565
rect -6913 -2615 -6793 -2599
rect -6735 -2565 -6615 -2518
rect -6735 -2599 -6719 -2565
rect -6631 -2599 -6615 -2565
rect -6735 -2615 -6615 -2599
rect -6557 -2565 -6437 -2518
rect -6557 -2599 -6541 -2565
rect -6453 -2599 -6437 -2565
rect -6557 -2615 -6437 -2599
rect -6379 -2565 -6259 -2518
rect -6379 -2599 -6363 -2565
rect -6275 -2599 -6259 -2565
rect -6379 -2615 -6259 -2599
rect -6201 -2565 -6081 -2518
rect -6201 -2599 -6185 -2565
rect -6097 -2599 -6081 -2565
rect -6201 -2615 -6081 -2599
rect -6023 -2565 -5903 -2518
rect -6023 -2599 -6007 -2565
rect -5919 -2599 -5903 -2565
rect -6023 -2615 -5903 -2599
rect -5845 -2565 -5725 -2518
rect -5845 -2599 -5829 -2565
rect -5741 -2599 -5725 -2565
rect -5845 -2615 -5725 -2599
rect -5667 -2565 -5547 -2518
rect -5667 -2599 -5651 -2565
rect -5563 -2599 -5547 -2565
rect -5667 -2615 -5547 -2599
rect -5489 -2565 -5369 -2518
rect -5489 -2599 -5473 -2565
rect -5385 -2599 -5369 -2565
rect -5489 -2615 -5369 -2599
rect -5311 -2565 -5191 -2518
rect -5311 -2599 -5295 -2565
rect -5207 -2599 -5191 -2565
rect -5311 -2615 -5191 -2599
rect -5133 -2565 -5013 -2518
rect -5133 -2599 -5117 -2565
rect -5029 -2599 -5013 -2565
rect -5133 -2615 -5013 -2599
rect -4955 -2565 -4835 -2518
rect -4955 -2599 -4939 -2565
rect -4851 -2599 -4835 -2565
rect -4955 -2615 -4835 -2599
rect -4777 -2565 -4657 -2518
rect -4777 -2599 -4761 -2565
rect -4673 -2599 -4657 -2565
rect -4777 -2615 -4657 -2599
rect -4599 -2565 -4479 -2518
rect -4599 -2599 -4583 -2565
rect -4495 -2599 -4479 -2565
rect -4599 -2615 -4479 -2599
rect -4421 -2565 -4301 -2518
rect -4421 -2599 -4405 -2565
rect -4317 -2599 -4301 -2565
rect -4421 -2615 -4301 -2599
rect -4243 -2565 -4123 -2518
rect -4243 -2599 -4227 -2565
rect -4139 -2599 -4123 -2565
rect -4243 -2615 -4123 -2599
rect -4065 -2565 -3945 -2518
rect -4065 -2599 -4049 -2565
rect -3961 -2599 -3945 -2565
rect -4065 -2615 -3945 -2599
rect -3887 -2565 -3767 -2518
rect -3887 -2599 -3871 -2565
rect -3783 -2599 -3767 -2565
rect -3887 -2615 -3767 -2599
rect -3709 -2565 -3589 -2518
rect -3709 -2599 -3693 -2565
rect -3605 -2599 -3589 -2565
rect -3709 -2615 -3589 -2599
rect -3531 -2565 -3411 -2518
rect -3531 -2599 -3515 -2565
rect -3427 -2599 -3411 -2565
rect -3531 -2615 -3411 -2599
rect -3353 -2565 -3233 -2518
rect -3353 -2599 -3337 -2565
rect -3249 -2599 -3233 -2565
rect -3353 -2615 -3233 -2599
rect -3175 -2565 -3055 -2518
rect -3175 -2599 -3159 -2565
rect -3071 -2599 -3055 -2565
rect -3175 -2615 -3055 -2599
rect -2997 -2565 -2877 -2518
rect -2997 -2599 -2981 -2565
rect -2893 -2599 -2877 -2565
rect -2997 -2615 -2877 -2599
rect -2819 -2565 -2699 -2518
rect -2819 -2599 -2803 -2565
rect -2715 -2599 -2699 -2565
rect -2819 -2615 -2699 -2599
rect -2641 -2565 -2521 -2518
rect -2641 -2599 -2625 -2565
rect -2537 -2599 -2521 -2565
rect -2641 -2615 -2521 -2599
rect -2463 -2565 -2343 -2518
rect -2463 -2599 -2447 -2565
rect -2359 -2599 -2343 -2565
rect -2463 -2615 -2343 -2599
rect -2285 -2565 -2165 -2518
rect -2285 -2599 -2269 -2565
rect -2181 -2599 -2165 -2565
rect -2285 -2615 -2165 -2599
rect -2107 -2565 -1987 -2518
rect -2107 -2599 -2091 -2565
rect -2003 -2599 -1987 -2565
rect -2107 -2615 -1987 -2599
rect -1929 -2565 -1809 -2518
rect -1929 -2599 -1913 -2565
rect -1825 -2599 -1809 -2565
rect -1929 -2615 -1809 -2599
rect -1751 -2565 -1631 -2518
rect -1751 -2599 -1735 -2565
rect -1647 -2599 -1631 -2565
rect -1751 -2615 -1631 -2599
rect -1573 -2565 -1453 -2518
rect -1573 -2599 -1557 -2565
rect -1469 -2599 -1453 -2565
rect -1573 -2615 -1453 -2599
rect -1395 -2565 -1275 -2518
rect -1395 -2599 -1379 -2565
rect -1291 -2599 -1275 -2565
rect -1395 -2615 -1275 -2599
rect -1217 -2565 -1097 -2518
rect -1217 -2599 -1201 -2565
rect -1113 -2599 -1097 -2565
rect -1217 -2615 -1097 -2599
rect -1039 -2565 -919 -2518
rect -1039 -2599 -1023 -2565
rect -935 -2599 -919 -2565
rect -1039 -2615 -919 -2599
rect -861 -2565 -741 -2518
rect -861 -2599 -845 -2565
rect -757 -2599 -741 -2565
rect -861 -2615 -741 -2599
rect -683 -2565 -563 -2518
rect -683 -2599 -667 -2565
rect -579 -2599 -563 -2565
rect -683 -2615 -563 -2599
rect -505 -2565 -385 -2518
rect -505 -2599 -489 -2565
rect -401 -2599 -385 -2565
rect -505 -2615 -385 -2599
rect -327 -2565 -207 -2518
rect -327 -2599 -311 -2565
rect -223 -2599 -207 -2565
rect -327 -2615 -207 -2599
rect -149 -2565 -29 -2518
rect -149 -2599 -133 -2565
rect -45 -2599 -29 -2565
rect -149 -2615 -29 -2599
rect 29 -2565 149 -2518
rect 29 -2599 45 -2565
rect 133 -2599 149 -2565
rect 29 -2615 149 -2599
rect 207 -2565 327 -2518
rect 207 -2599 223 -2565
rect 311 -2599 327 -2565
rect 207 -2615 327 -2599
rect 385 -2565 505 -2518
rect 385 -2599 401 -2565
rect 489 -2599 505 -2565
rect 385 -2615 505 -2599
rect 563 -2565 683 -2518
rect 563 -2599 579 -2565
rect 667 -2599 683 -2565
rect 563 -2615 683 -2599
rect 741 -2565 861 -2518
rect 741 -2599 757 -2565
rect 845 -2599 861 -2565
rect 741 -2615 861 -2599
rect 919 -2565 1039 -2518
rect 919 -2599 935 -2565
rect 1023 -2599 1039 -2565
rect 919 -2615 1039 -2599
rect 1097 -2565 1217 -2518
rect 1097 -2599 1113 -2565
rect 1201 -2599 1217 -2565
rect 1097 -2615 1217 -2599
rect 1275 -2565 1395 -2518
rect 1275 -2599 1291 -2565
rect 1379 -2599 1395 -2565
rect 1275 -2615 1395 -2599
rect 1453 -2565 1573 -2518
rect 1453 -2599 1469 -2565
rect 1557 -2599 1573 -2565
rect 1453 -2615 1573 -2599
rect 1631 -2565 1751 -2518
rect 1631 -2599 1647 -2565
rect 1735 -2599 1751 -2565
rect 1631 -2615 1751 -2599
rect 1809 -2565 1929 -2518
rect 1809 -2599 1825 -2565
rect 1913 -2599 1929 -2565
rect 1809 -2615 1929 -2599
rect 1987 -2565 2107 -2518
rect 1987 -2599 2003 -2565
rect 2091 -2599 2107 -2565
rect 1987 -2615 2107 -2599
rect 2165 -2565 2285 -2518
rect 2165 -2599 2181 -2565
rect 2269 -2599 2285 -2565
rect 2165 -2615 2285 -2599
rect 2343 -2565 2463 -2518
rect 2343 -2599 2359 -2565
rect 2447 -2599 2463 -2565
rect 2343 -2615 2463 -2599
rect 2521 -2565 2641 -2518
rect 2521 -2599 2537 -2565
rect 2625 -2599 2641 -2565
rect 2521 -2615 2641 -2599
rect 2699 -2565 2819 -2518
rect 2699 -2599 2715 -2565
rect 2803 -2599 2819 -2565
rect 2699 -2615 2819 -2599
rect 2877 -2565 2997 -2518
rect 2877 -2599 2893 -2565
rect 2981 -2599 2997 -2565
rect 2877 -2615 2997 -2599
rect 3055 -2565 3175 -2518
rect 3055 -2599 3071 -2565
rect 3159 -2599 3175 -2565
rect 3055 -2615 3175 -2599
rect 3233 -2565 3353 -2518
rect 3233 -2599 3249 -2565
rect 3337 -2599 3353 -2565
rect 3233 -2615 3353 -2599
rect 3411 -2565 3531 -2518
rect 3411 -2599 3427 -2565
rect 3515 -2599 3531 -2565
rect 3411 -2615 3531 -2599
rect 3589 -2565 3709 -2518
rect 3589 -2599 3605 -2565
rect 3693 -2599 3709 -2565
rect 3589 -2615 3709 -2599
rect 3767 -2565 3887 -2518
rect 3767 -2599 3783 -2565
rect 3871 -2599 3887 -2565
rect 3767 -2615 3887 -2599
rect 3945 -2565 4065 -2518
rect 3945 -2599 3961 -2565
rect 4049 -2599 4065 -2565
rect 3945 -2615 4065 -2599
rect 4123 -2565 4243 -2518
rect 4123 -2599 4139 -2565
rect 4227 -2599 4243 -2565
rect 4123 -2615 4243 -2599
rect 4301 -2565 4421 -2518
rect 4301 -2599 4317 -2565
rect 4405 -2599 4421 -2565
rect 4301 -2615 4421 -2599
rect 4479 -2565 4599 -2518
rect 4479 -2599 4495 -2565
rect 4583 -2599 4599 -2565
rect 4479 -2615 4599 -2599
rect 4657 -2565 4777 -2518
rect 4657 -2599 4673 -2565
rect 4761 -2599 4777 -2565
rect 4657 -2615 4777 -2599
rect 4835 -2565 4955 -2518
rect 4835 -2599 4851 -2565
rect 4939 -2599 4955 -2565
rect 4835 -2615 4955 -2599
rect 5013 -2565 5133 -2518
rect 5013 -2599 5029 -2565
rect 5117 -2599 5133 -2565
rect 5013 -2615 5133 -2599
rect 5191 -2565 5311 -2518
rect 5191 -2599 5207 -2565
rect 5295 -2599 5311 -2565
rect 5191 -2615 5311 -2599
rect 5369 -2565 5489 -2518
rect 5369 -2599 5385 -2565
rect 5473 -2599 5489 -2565
rect 5369 -2615 5489 -2599
rect 5547 -2565 5667 -2518
rect 5547 -2599 5563 -2565
rect 5651 -2599 5667 -2565
rect 5547 -2615 5667 -2599
rect 5725 -2565 5845 -2518
rect 5725 -2599 5741 -2565
rect 5829 -2599 5845 -2565
rect 5725 -2615 5845 -2599
rect 5903 -2565 6023 -2518
rect 5903 -2599 5919 -2565
rect 6007 -2599 6023 -2565
rect 5903 -2615 6023 -2599
rect 6081 -2565 6201 -2518
rect 6081 -2599 6097 -2565
rect 6185 -2599 6201 -2565
rect 6081 -2615 6201 -2599
rect 6259 -2565 6379 -2518
rect 6259 -2599 6275 -2565
rect 6363 -2599 6379 -2565
rect 6259 -2615 6379 -2599
rect 6437 -2565 6557 -2518
rect 6437 -2599 6453 -2565
rect 6541 -2599 6557 -2565
rect 6437 -2615 6557 -2599
rect 6615 -2565 6735 -2518
rect 6615 -2599 6631 -2565
rect 6719 -2599 6735 -2565
rect 6615 -2615 6735 -2599
rect 6793 -2565 6913 -2518
rect 6793 -2599 6809 -2565
rect 6897 -2599 6913 -2565
rect 6793 -2615 6913 -2599
rect 6971 -2565 7091 -2518
rect 6971 -2599 6987 -2565
rect 7075 -2599 7091 -2565
rect 6971 -2615 7091 -2599
rect 7149 -2565 7269 -2518
rect 7149 -2599 7165 -2565
rect 7253 -2599 7269 -2565
rect 7149 -2615 7269 -2599
rect 7327 -2565 7447 -2518
rect 7327 -2599 7343 -2565
rect 7431 -2599 7447 -2565
rect 7327 -2615 7447 -2599
rect 7505 -2565 7625 -2518
rect 7505 -2599 7521 -2565
rect 7609 -2599 7625 -2565
rect 7505 -2615 7625 -2599
rect 7683 -2565 7803 -2518
rect 7683 -2599 7699 -2565
rect 7787 -2599 7803 -2565
rect 7683 -2615 7803 -2599
rect 7861 -2565 7981 -2518
rect 7861 -2599 7877 -2565
rect 7965 -2599 7981 -2565
rect 7861 -2615 7981 -2599
rect 8039 -2565 8159 -2518
rect 8039 -2599 8055 -2565
rect 8143 -2599 8159 -2565
rect 8039 -2615 8159 -2599
rect 8217 -2565 8337 -2518
rect 8217 -2599 8233 -2565
rect 8321 -2599 8337 -2565
rect 8217 -2615 8337 -2599
rect 8395 -2565 8515 -2518
rect 8395 -2599 8411 -2565
rect 8499 -2599 8515 -2565
rect 8395 -2615 8515 -2599
rect 8573 -2565 8693 -2518
rect 8573 -2599 8589 -2565
rect 8677 -2599 8693 -2565
rect 8573 -2615 8693 -2599
rect 8751 -2565 8871 -2518
rect 8751 -2599 8767 -2565
rect 8855 -2599 8871 -2565
rect 8751 -2615 8871 -2599
<< polycont >>
rect -8855 2565 -8767 2599
rect -8677 2565 -8589 2599
rect -8499 2565 -8411 2599
rect -8321 2565 -8233 2599
rect -8143 2565 -8055 2599
rect -7965 2565 -7877 2599
rect -7787 2565 -7699 2599
rect -7609 2565 -7521 2599
rect -7431 2565 -7343 2599
rect -7253 2565 -7165 2599
rect -7075 2565 -6987 2599
rect -6897 2565 -6809 2599
rect -6719 2565 -6631 2599
rect -6541 2565 -6453 2599
rect -6363 2565 -6275 2599
rect -6185 2565 -6097 2599
rect -6007 2565 -5919 2599
rect -5829 2565 -5741 2599
rect -5651 2565 -5563 2599
rect -5473 2565 -5385 2599
rect -5295 2565 -5207 2599
rect -5117 2565 -5029 2599
rect -4939 2565 -4851 2599
rect -4761 2565 -4673 2599
rect -4583 2565 -4495 2599
rect -4405 2565 -4317 2599
rect -4227 2565 -4139 2599
rect -4049 2565 -3961 2599
rect -3871 2565 -3783 2599
rect -3693 2565 -3605 2599
rect -3515 2565 -3427 2599
rect -3337 2565 -3249 2599
rect -3159 2565 -3071 2599
rect -2981 2565 -2893 2599
rect -2803 2565 -2715 2599
rect -2625 2565 -2537 2599
rect -2447 2565 -2359 2599
rect -2269 2565 -2181 2599
rect -2091 2565 -2003 2599
rect -1913 2565 -1825 2599
rect -1735 2565 -1647 2599
rect -1557 2565 -1469 2599
rect -1379 2565 -1291 2599
rect -1201 2565 -1113 2599
rect -1023 2565 -935 2599
rect -845 2565 -757 2599
rect -667 2565 -579 2599
rect -489 2565 -401 2599
rect -311 2565 -223 2599
rect -133 2565 -45 2599
rect 45 2565 133 2599
rect 223 2565 311 2599
rect 401 2565 489 2599
rect 579 2565 667 2599
rect 757 2565 845 2599
rect 935 2565 1023 2599
rect 1113 2565 1201 2599
rect 1291 2565 1379 2599
rect 1469 2565 1557 2599
rect 1647 2565 1735 2599
rect 1825 2565 1913 2599
rect 2003 2565 2091 2599
rect 2181 2565 2269 2599
rect 2359 2565 2447 2599
rect 2537 2565 2625 2599
rect 2715 2565 2803 2599
rect 2893 2565 2981 2599
rect 3071 2565 3159 2599
rect 3249 2565 3337 2599
rect 3427 2565 3515 2599
rect 3605 2565 3693 2599
rect 3783 2565 3871 2599
rect 3961 2565 4049 2599
rect 4139 2565 4227 2599
rect 4317 2565 4405 2599
rect 4495 2565 4583 2599
rect 4673 2565 4761 2599
rect 4851 2565 4939 2599
rect 5029 2565 5117 2599
rect 5207 2565 5295 2599
rect 5385 2565 5473 2599
rect 5563 2565 5651 2599
rect 5741 2565 5829 2599
rect 5919 2565 6007 2599
rect 6097 2565 6185 2599
rect 6275 2565 6363 2599
rect 6453 2565 6541 2599
rect 6631 2565 6719 2599
rect 6809 2565 6897 2599
rect 6987 2565 7075 2599
rect 7165 2565 7253 2599
rect 7343 2565 7431 2599
rect 7521 2565 7609 2599
rect 7699 2565 7787 2599
rect 7877 2565 7965 2599
rect 8055 2565 8143 2599
rect 8233 2565 8321 2599
rect 8411 2565 8499 2599
rect 8589 2565 8677 2599
rect 8767 2565 8855 2599
rect -8855 37 -8767 71
rect -8677 37 -8589 71
rect -8499 37 -8411 71
rect -8321 37 -8233 71
rect -8143 37 -8055 71
rect -7965 37 -7877 71
rect -7787 37 -7699 71
rect -7609 37 -7521 71
rect -7431 37 -7343 71
rect -7253 37 -7165 71
rect -7075 37 -6987 71
rect -6897 37 -6809 71
rect -6719 37 -6631 71
rect -6541 37 -6453 71
rect -6363 37 -6275 71
rect -6185 37 -6097 71
rect -6007 37 -5919 71
rect -5829 37 -5741 71
rect -5651 37 -5563 71
rect -5473 37 -5385 71
rect -5295 37 -5207 71
rect -5117 37 -5029 71
rect -4939 37 -4851 71
rect -4761 37 -4673 71
rect -4583 37 -4495 71
rect -4405 37 -4317 71
rect -4227 37 -4139 71
rect -4049 37 -3961 71
rect -3871 37 -3783 71
rect -3693 37 -3605 71
rect -3515 37 -3427 71
rect -3337 37 -3249 71
rect -3159 37 -3071 71
rect -2981 37 -2893 71
rect -2803 37 -2715 71
rect -2625 37 -2537 71
rect -2447 37 -2359 71
rect -2269 37 -2181 71
rect -2091 37 -2003 71
rect -1913 37 -1825 71
rect -1735 37 -1647 71
rect -1557 37 -1469 71
rect -1379 37 -1291 71
rect -1201 37 -1113 71
rect -1023 37 -935 71
rect -845 37 -757 71
rect -667 37 -579 71
rect -489 37 -401 71
rect -311 37 -223 71
rect -133 37 -45 71
rect 45 37 133 71
rect 223 37 311 71
rect 401 37 489 71
rect 579 37 667 71
rect 757 37 845 71
rect 935 37 1023 71
rect 1113 37 1201 71
rect 1291 37 1379 71
rect 1469 37 1557 71
rect 1647 37 1735 71
rect 1825 37 1913 71
rect 2003 37 2091 71
rect 2181 37 2269 71
rect 2359 37 2447 71
rect 2537 37 2625 71
rect 2715 37 2803 71
rect 2893 37 2981 71
rect 3071 37 3159 71
rect 3249 37 3337 71
rect 3427 37 3515 71
rect 3605 37 3693 71
rect 3783 37 3871 71
rect 3961 37 4049 71
rect 4139 37 4227 71
rect 4317 37 4405 71
rect 4495 37 4583 71
rect 4673 37 4761 71
rect 4851 37 4939 71
rect 5029 37 5117 71
rect 5207 37 5295 71
rect 5385 37 5473 71
rect 5563 37 5651 71
rect 5741 37 5829 71
rect 5919 37 6007 71
rect 6097 37 6185 71
rect 6275 37 6363 71
rect 6453 37 6541 71
rect 6631 37 6719 71
rect 6809 37 6897 71
rect 6987 37 7075 71
rect 7165 37 7253 71
rect 7343 37 7431 71
rect 7521 37 7609 71
rect 7699 37 7787 71
rect 7877 37 7965 71
rect 8055 37 8143 71
rect 8233 37 8321 71
rect 8411 37 8499 71
rect 8589 37 8677 71
rect 8767 37 8855 71
rect -8855 -71 -8767 -37
rect -8677 -71 -8589 -37
rect -8499 -71 -8411 -37
rect -8321 -71 -8233 -37
rect -8143 -71 -8055 -37
rect -7965 -71 -7877 -37
rect -7787 -71 -7699 -37
rect -7609 -71 -7521 -37
rect -7431 -71 -7343 -37
rect -7253 -71 -7165 -37
rect -7075 -71 -6987 -37
rect -6897 -71 -6809 -37
rect -6719 -71 -6631 -37
rect -6541 -71 -6453 -37
rect -6363 -71 -6275 -37
rect -6185 -71 -6097 -37
rect -6007 -71 -5919 -37
rect -5829 -71 -5741 -37
rect -5651 -71 -5563 -37
rect -5473 -71 -5385 -37
rect -5295 -71 -5207 -37
rect -5117 -71 -5029 -37
rect -4939 -71 -4851 -37
rect -4761 -71 -4673 -37
rect -4583 -71 -4495 -37
rect -4405 -71 -4317 -37
rect -4227 -71 -4139 -37
rect -4049 -71 -3961 -37
rect -3871 -71 -3783 -37
rect -3693 -71 -3605 -37
rect -3515 -71 -3427 -37
rect -3337 -71 -3249 -37
rect -3159 -71 -3071 -37
rect -2981 -71 -2893 -37
rect -2803 -71 -2715 -37
rect -2625 -71 -2537 -37
rect -2447 -71 -2359 -37
rect -2269 -71 -2181 -37
rect -2091 -71 -2003 -37
rect -1913 -71 -1825 -37
rect -1735 -71 -1647 -37
rect -1557 -71 -1469 -37
rect -1379 -71 -1291 -37
rect -1201 -71 -1113 -37
rect -1023 -71 -935 -37
rect -845 -71 -757 -37
rect -667 -71 -579 -37
rect -489 -71 -401 -37
rect -311 -71 -223 -37
rect -133 -71 -45 -37
rect 45 -71 133 -37
rect 223 -71 311 -37
rect 401 -71 489 -37
rect 579 -71 667 -37
rect 757 -71 845 -37
rect 935 -71 1023 -37
rect 1113 -71 1201 -37
rect 1291 -71 1379 -37
rect 1469 -71 1557 -37
rect 1647 -71 1735 -37
rect 1825 -71 1913 -37
rect 2003 -71 2091 -37
rect 2181 -71 2269 -37
rect 2359 -71 2447 -37
rect 2537 -71 2625 -37
rect 2715 -71 2803 -37
rect 2893 -71 2981 -37
rect 3071 -71 3159 -37
rect 3249 -71 3337 -37
rect 3427 -71 3515 -37
rect 3605 -71 3693 -37
rect 3783 -71 3871 -37
rect 3961 -71 4049 -37
rect 4139 -71 4227 -37
rect 4317 -71 4405 -37
rect 4495 -71 4583 -37
rect 4673 -71 4761 -37
rect 4851 -71 4939 -37
rect 5029 -71 5117 -37
rect 5207 -71 5295 -37
rect 5385 -71 5473 -37
rect 5563 -71 5651 -37
rect 5741 -71 5829 -37
rect 5919 -71 6007 -37
rect 6097 -71 6185 -37
rect 6275 -71 6363 -37
rect 6453 -71 6541 -37
rect 6631 -71 6719 -37
rect 6809 -71 6897 -37
rect 6987 -71 7075 -37
rect 7165 -71 7253 -37
rect 7343 -71 7431 -37
rect 7521 -71 7609 -37
rect 7699 -71 7787 -37
rect 7877 -71 7965 -37
rect 8055 -71 8143 -37
rect 8233 -71 8321 -37
rect 8411 -71 8499 -37
rect 8589 -71 8677 -37
rect 8767 -71 8855 -37
rect -8855 -2599 -8767 -2565
rect -8677 -2599 -8589 -2565
rect -8499 -2599 -8411 -2565
rect -8321 -2599 -8233 -2565
rect -8143 -2599 -8055 -2565
rect -7965 -2599 -7877 -2565
rect -7787 -2599 -7699 -2565
rect -7609 -2599 -7521 -2565
rect -7431 -2599 -7343 -2565
rect -7253 -2599 -7165 -2565
rect -7075 -2599 -6987 -2565
rect -6897 -2599 -6809 -2565
rect -6719 -2599 -6631 -2565
rect -6541 -2599 -6453 -2565
rect -6363 -2599 -6275 -2565
rect -6185 -2599 -6097 -2565
rect -6007 -2599 -5919 -2565
rect -5829 -2599 -5741 -2565
rect -5651 -2599 -5563 -2565
rect -5473 -2599 -5385 -2565
rect -5295 -2599 -5207 -2565
rect -5117 -2599 -5029 -2565
rect -4939 -2599 -4851 -2565
rect -4761 -2599 -4673 -2565
rect -4583 -2599 -4495 -2565
rect -4405 -2599 -4317 -2565
rect -4227 -2599 -4139 -2565
rect -4049 -2599 -3961 -2565
rect -3871 -2599 -3783 -2565
rect -3693 -2599 -3605 -2565
rect -3515 -2599 -3427 -2565
rect -3337 -2599 -3249 -2565
rect -3159 -2599 -3071 -2565
rect -2981 -2599 -2893 -2565
rect -2803 -2599 -2715 -2565
rect -2625 -2599 -2537 -2565
rect -2447 -2599 -2359 -2565
rect -2269 -2599 -2181 -2565
rect -2091 -2599 -2003 -2565
rect -1913 -2599 -1825 -2565
rect -1735 -2599 -1647 -2565
rect -1557 -2599 -1469 -2565
rect -1379 -2599 -1291 -2565
rect -1201 -2599 -1113 -2565
rect -1023 -2599 -935 -2565
rect -845 -2599 -757 -2565
rect -667 -2599 -579 -2565
rect -489 -2599 -401 -2565
rect -311 -2599 -223 -2565
rect -133 -2599 -45 -2565
rect 45 -2599 133 -2565
rect 223 -2599 311 -2565
rect 401 -2599 489 -2565
rect 579 -2599 667 -2565
rect 757 -2599 845 -2565
rect 935 -2599 1023 -2565
rect 1113 -2599 1201 -2565
rect 1291 -2599 1379 -2565
rect 1469 -2599 1557 -2565
rect 1647 -2599 1735 -2565
rect 1825 -2599 1913 -2565
rect 2003 -2599 2091 -2565
rect 2181 -2599 2269 -2565
rect 2359 -2599 2447 -2565
rect 2537 -2599 2625 -2565
rect 2715 -2599 2803 -2565
rect 2893 -2599 2981 -2565
rect 3071 -2599 3159 -2565
rect 3249 -2599 3337 -2565
rect 3427 -2599 3515 -2565
rect 3605 -2599 3693 -2565
rect 3783 -2599 3871 -2565
rect 3961 -2599 4049 -2565
rect 4139 -2599 4227 -2565
rect 4317 -2599 4405 -2565
rect 4495 -2599 4583 -2565
rect 4673 -2599 4761 -2565
rect 4851 -2599 4939 -2565
rect 5029 -2599 5117 -2565
rect 5207 -2599 5295 -2565
rect 5385 -2599 5473 -2565
rect 5563 -2599 5651 -2565
rect 5741 -2599 5829 -2565
rect 5919 -2599 6007 -2565
rect 6097 -2599 6185 -2565
rect 6275 -2599 6363 -2565
rect 6453 -2599 6541 -2565
rect 6631 -2599 6719 -2565
rect 6809 -2599 6897 -2565
rect 6987 -2599 7075 -2565
rect 7165 -2599 7253 -2565
rect 7343 -2599 7431 -2565
rect 7521 -2599 7609 -2565
rect 7699 -2599 7787 -2565
rect 7877 -2599 7965 -2565
rect 8055 -2599 8143 -2565
rect 8233 -2599 8321 -2565
rect 8411 -2599 8499 -2565
rect 8589 -2599 8677 -2565
rect 8767 -2599 8855 -2565
<< locali >>
rect -9031 2667 -8935 2701
rect 8935 2667 9031 2701
rect -9031 2605 -8997 2667
rect 8997 2605 9031 2667
rect -8871 2565 -8855 2599
rect -8767 2565 -8751 2599
rect -8693 2565 -8677 2599
rect -8589 2565 -8573 2599
rect -8515 2565 -8499 2599
rect -8411 2565 -8395 2599
rect -8337 2565 -8321 2599
rect -8233 2565 -8217 2599
rect -8159 2565 -8143 2599
rect -8055 2565 -8039 2599
rect -7981 2565 -7965 2599
rect -7877 2565 -7861 2599
rect -7803 2565 -7787 2599
rect -7699 2565 -7683 2599
rect -7625 2565 -7609 2599
rect -7521 2565 -7505 2599
rect -7447 2565 -7431 2599
rect -7343 2565 -7327 2599
rect -7269 2565 -7253 2599
rect -7165 2565 -7149 2599
rect -7091 2565 -7075 2599
rect -6987 2565 -6971 2599
rect -6913 2565 -6897 2599
rect -6809 2565 -6793 2599
rect -6735 2565 -6719 2599
rect -6631 2565 -6615 2599
rect -6557 2565 -6541 2599
rect -6453 2565 -6437 2599
rect -6379 2565 -6363 2599
rect -6275 2565 -6259 2599
rect -6201 2565 -6185 2599
rect -6097 2565 -6081 2599
rect -6023 2565 -6007 2599
rect -5919 2565 -5903 2599
rect -5845 2565 -5829 2599
rect -5741 2565 -5725 2599
rect -5667 2565 -5651 2599
rect -5563 2565 -5547 2599
rect -5489 2565 -5473 2599
rect -5385 2565 -5369 2599
rect -5311 2565 -5295 2599
rect -5207 2565 -5191 2599
rect -5133 2565 -5117 2599
rect -5029 2565 -5013 2599
rect -4955 2565 -4939 2599
rect -4851 2565 -4835 2599
rect -4777 2565 -4761 2599
rect -4673 2565 -4657 2599
rect -4599 2565 -4583 2599
rect -4495 2565 -4479 2599
rect -4421 2565 -4405 2599
rect -4317 2565 -4301 2599
rect -4243 2565 -4227 2599
rect -4139 2565 -4123 2599
rect -4065 2565 -4049 2599
rect -3961 2565 -3945 2599
rect -3887 2565 -3871 2599
rect -3783 2565 -3767 2599
rect -3709 2565 -3693 2599
rect -3605 2565 -3589 2599
rect -3531 2565 -3515 2599
rect -3427 2565 -3411 2599
rect -3353 2565 -3337 2599
rect -3249 2565 -3233 2599
rect -3175 2565 -3159 2599
rect -3071 2565 -3055 2599
rect -2997 2565 -2981 2599
rect -2893 2565 -2877 2599
rect -2819 2565 -2803 2599
rect -2715 2565 -2699 2599
rect -2641 2565 -2625 2599
rect -2537 2565 -2521 2599
rect -2463 2565 -2447 2599
rect -2359 2565 -2343 2599
rect -2285 2565 -2269 2599
rect -2181 2565 -2165 2599
rect -2107 2565 -2091 2599
rect -2003 2565 -1987 2599
rect -1929 2565 -1913 2599
rect -1825 2565 -1809 2599
rect -1751 2565 -1735 2599
rect -1647 2565 -1631 2599
rect -1573 2565 -1557 2599
rect -1469 2565 -1453 2599
rect -1395 2565 -1379 2599
rect -1291 2565 -1275 2599
rect -1217 2565 -1201 2599
rect -1113 2565 -1097 2599
rect -1039 2565 -1023 2599
rect -935 2565 -919 2599
rect -861 2565 -845 2599
rect -757 2565 -741 2599
rect -683 2565 -667 2599
rect -579 2565 -563 2599
rect -505 2565 -489 2599
rect -401 2565 -385 2599
rect -327 2565 -311 2599
rect -223 2565 -207 2599
rect -149 2565 -133 2599
rect -45 2565 -29 2599
rect 29 2565 45 2599
rect 133 2565 149 2599
rect 207 2565 223 2599
rect 311 2565 327 2599
rect 385 2565 401 2599
rect 489 2565 505 2599
rect 563 2565 579 2599
rect 667 2565 683 2599
rect 741 2565 757 2599
rect 845 2565 861 2599
rect 919 2565 935 2599
rect 1023 2565 1039 2599
rect 1097 2565 1113 2599
rect 1201 2565 1217 2599
rect 1275 2565 1291 2599
rect 1379 2565 1395 2599
rect 1453 2565 1469 2599
rect 1557 2565 1573 2599
rect 1631 2565 1647 2599
rect 1735 2565 1751 2599
rect 1809 2565 1825 2599
rect 1913 2565 1929 2599
rect 1987 2565 2003 2599
rect 2091 2565 2107 2599
rect 2165 2565 2181 2599
rect 2269 2565 2285 2599
rect 2343 2565 2359 2599
rect 2447 2565 2463 2599
rect 2521 2565 2537 2599
rect 2625 2565 2641 2599
rect 2699 2565 2715 2599
rect 2803 2565 2819 2599
rect 2877 2565 2893 2599
rect 2981 2565 2997 2599
rect 3055 2565 3071 2599
rect 3159 2565 3175 2599
rect 3233 2565 3249 2599
rect 3337 2565 3353 2599
rect 3411 2565 3427 2599
rect 3515 2565 3531 2599
rect 3589 2565 3605 2599
rect 3693 2565 3709 2599
rect 3767 2565 3783 2599
rect 3871 2565 3887 2599
rect 3945 2565 3961 2599
rect 4049 2565 4065 2599
rect 4123 2565 4139 2599
rect 4227 2565 4243 2599
rect 4301 2565 4317 2599
rect 4405 2565 4421 2599
rect 4479 2565 4495 2599
rect 4583 2565 4599 2599
rect 4657 2565 4673 2599
rect 4761 2565 4777 2599
rect 4835 2565 4851 2599
rect 4939 2565 4955 2599
rect 5013 2565 5029 2599
rect 5117 2565 5133 2599
rect 5191 2565 5207 2599
rect 5295 2565 5311 2599
rect 5369 2565 5385 2599
rect 5473 2565 5489 2599
rect 5547 2565 5563 2599
rect 5651 2565 5667 2599
rect 5725 2565 5741 2599
rect 5829 2565 5845 2599
rect 5903 2565 5919 2599
rect 6007 2565 6023 2599
rect 6081 2565 6097 2599
rect 6185 2565 6201 2599
rect 6259 2565 6275 2599
rect 6363 2565 6379 2599
rect 6437 2565 6453 2599
rect 6541 2565 6557 2599
rect 6615 2565 6631 2599
rect 6719 2565 6735 2599
rect 6793 2565 6809 2599
rect 6897 2565 6913 2599
rect 6971 2565 6987 2599
rect 7075 2565 7091 2599
rect 7149 2565 7165 2599
rect 7253 2565 7269 2599
rect 7327 2565 7343 2599
rect 7431 2565 7447 2599
rect 7505 2565 7521 2599
rect 7609 2565 7625 2599
rect 7683 2565 7699 2599
rect 7787 2565 7803 2599
rect 7861 2565 7877 2599
rect 7965 2565 7981 2599
rect 8039 2565 8055 2599
rect 8143 2565 8159 2599
rect 8217 2565 8233 2599
rect 8321 2565 8337 2599
rect 8395 2565 8411 2599
rect 8499 2565 8515 2599
rect 8573 2565 8589 2599
rect 8677 2565 8693 2599
rect 8751 2565 8767 2599
rect 8855 2565 8871 2599
rect -8917 2506 -8883 2522
rect -8917 114 -8883 130
rect -8739 2506 -8705 2522
rect -8739 114 -8705 130
rect -8561 2506 -8527 2522
rect -8561 114 -8527 130
rect -8383 2506 -8349 2522
rect -8383 114 -8349 130
rect -8205 2506 -8171 2522
rect -8205 114 -8171 130
rect -8027 2506 -7993 2522
rect -8027 114 -7993 130
rect -7849 2506 -7815 2522
rect -7849 114 -7815 130
rect -7671 2506 -7637 2522
rect -7671 114 -7637 130
rect -7493 2506 -7459 2522
rect -7493 114 -7459 130
rect -7315 2506 -7281 2522
rect -7315 114 -7281 130
rect -7137 2506 -7103 2522
rect -7137 114 -7103 130
rect -6959 2506 -6925 2522
rect -6959 114 -6925 130
rect -6781 2506 -6747 2522
rect -6781 114 -6747 130
rect -6603 2506 -6569 2522
rect -6603 114 -6569 130
rect -6425 2506 -6391 2522
rect -6425 114 -6391 130
rect -6247 2506 -6213 2522
rect -6247 114 -6213 130
rect -6069 2506 -6035 2522
rect -6069 114 -6035 130
rect -5891 2506 -5857 2522
rect -5891 114 -5857 130
rect -5713 2506 -5679 2522
rect -5713 114 -5679 130
rect -5535 2506 -5501 2522
rect -5535 114 -5501 130
rect -5357 2506 -5323 2522
rect -5357 114 -5323 130
rect -5179 2506 -5145 2522
rect -5179 114 -5145 130
rect -5001 2506 -4967 2522
rect -5001 114 -4967 130
rect -4823 2506 -4789 2522
rect -4823 114 -4789 130
rect -4645 2506 -4611 2522
rect -4645 114 -4611 130
rect -4467 2506 -4433 2522
rect -4467 114 -4433 130
rect -4289 2506 -4255 2522
rect -4289 114 -4255 130
rect -4111 2506 -4077 2522
rect -4111 114 -4077 130
rect -3933 2506 -3899 2522
rect -3933 114 -3899 130
rect -3755 2506 -3721 2522
rect -3755 114 -3721 130
rect -3577 2506 -3543 2522
rect -3577 114 -3543 130
rect -3399 2506 -3365 2522
rect -3399 114 -3365 130
rect -3221 2506 -3187 2522
rect -3221 114 -3187 130
rect -3043 2506 -3009 2522
rect -3043 114 -3009 130
rect -2865 2506 -2831 2522
rect -2865 114 -2831 130
rect -2687 2506 -2653 2522
rect -2687 114 -2653 130
rect -2509 2506 -2475 2522
rect -2509 114 -2475 130
rect -2331 2506 -2297 2522
rect -2331 114 -2297 130
rect -2153 2506 -2119 2522
rect -2153 114 -2119 130
rect -1975 2506 -1941 2522
rect -1975 114 -1941 130
rect -1797 2506 -1763 2522
rect -1797 114 -1763 130
rect -1619 2506 -1585 2522
rect -1619 114 -1585 130
rect -1441 2506 -1407 2522
rect -1441 114 -1407 130
rect -1263 2506 -1229 2522
rect -1263 114 -1229 130
rect -1085 2506 -1051 2522
rect -1085 114 -1051 130
rect -907 2506 -873 2522
rect -907 114 -873 130
rect -729 2506 -695 2522
rect -729 114 -695 130
rect -551 2506 -517 2522
rect -551 114 -517 130
rect -373 2506 -339 2522
rect -373 114 -339 130
rect -195 2506 -161 2522
rect -195 114 -161 130
rect -17 2506 17 2522
rect -17 114 17 130
rect 161 2506 195 2522
rect 161 114 195 130
rect 339 2506 373 2522
rect 339 114 373 130
rect 517 2506 551 2522
rect 517 114 551 130
rect 695 2506 729 2522
rect 695 114 729 130
rect 873 2506 907 2522
rect 873 114 907 130
rect 1051 2506 1085 2522
rect 1051 114 1085 130
rect 1229 2506 1263 2522
rect 1229 114 1263 130
rect 1407 2506 1441 2522
rect 1407 114 1441 130
rect 1585 2506 1619 2522
rect 1585 114 1619 130
rect 1763 2506 1797 2522
rect 1763 114 1797 130
rect 1941 2506 1975 2522
rect 1941 114 1975 130
rect 2119 2506 2153 2522
rect 2119 114 2153 130
rect 2297 2506 2331 2522
rect 2297 114 2331 130
rect 2475 2506 2509 2522
rect 2475 114 2509 130
rect 2653 2506 2687 2522
rect 2653 114 2687 130
rect 2831 2506 2865 2522
rect 2831 114 2865 130
rect 3009 2506 3043 2522
rect 3009 114 3043 130
rect 3187 2506 3221 2522
rect 3187 114 3221 130
rect 3365 2506 3399 2522
rect 3365 114 3399 130
rect 3543 2506 3577 2522
rect 3543 114 3577 130
rect 3721 2506 3755 2522
rect 3721 114 3755 130
rect 3899 2506 3933 2522
rect 3899 114 3933 130
rect 4077 2506 4111 2522
rect 4077 114 4111 130
rect 4255 2506 4289 2522
rect 4255 114 4289 130
rect 4433 2506 4467 2522
rect 4433 114 4467 130
rect 4611 2506 4645 2522
rect 4611 114 4645 130
rect 4789 2506 4823 2522
rect 4789 114 4823 130
rect 4967 2506 5001 2522
rect 4967 114 5001 130
rect 5145 2506 5179 2522
rect 5145 114 5179 130
rect 5323 2506 5357 2522
rect 5323 114 5357 130
rect 5501 2506 5535 2522
rect 5501 114 5535 130
rect 5679 2506 5713 2522
rect 5679 114 5713 130
rect 5857 2506 5891 2522
rect 5857 114 5891 130
rect 6035 2506 6069 2522
rect 6035 114 6069 130
rect 6213 2506 6247 2522
rect 6213 114 6247 130
rect 6391 2506 6425 2522
rect 6391 114 6425 130
rect 6569 2506 6603 2522
rect 6569 114 6603 130
rect 6747 2506 6781 2522
rect 6747 114 6781 130
rect 6925 2506 6959 2522
rect 6925 114 6959 130
rect 7103 2506 7137 2522
rect 7103 114 7137 130
rect 7281 2506 7315 2522
rect 7281 114 7315 130
rect 7459 2506 7493 2522
rect 7459 114 7493 130
rect 7637 2506 7671 2522
rect 7637 114 7671 130
rect 7815 2506 7849 2522
rect 7815 114 7849 130
rect 7993 2506 8027 2522
rect 7993 114 8027 130
rect 8171 2506 8205 2522
rect 8171 114 8205 130
rect 8349 2506 8383 2522
rect 8349 114 8383 130
rect 8527 2506 8561 2522
rect 8527 114 8561 130
rect 8705 2506 8739 2522
rect 8705 114 8739 130
rect 8883 2506 8917 2522
rect 8883 114 8917 130
rect -8871 37 -8855 71
rect -8767 37 -8751 71
rect -8693 37 -8677 71
rect -8589 37 -8573 71
rect -8515 37 -8499 71
rect -8411 37 -8395 71
rect -8337 37 -8321 71
rect -8233 37 -8217 71
rect -8159 37 -8143 71
rect -8055 37 -8039 71
rect -7981 37 -7965 71
rect -7877 37 -7861 71
rect -7803 37 -7787 71
rect -7699 37 -7683 71
rect -7625 37 -7609 71
rect -7521 37 -7505 71
rect -7447 37 -7431 71
rect -7343 37 -7327 71
rect -7269 37 -7253 71
rect -7165 37 -7149 71
rect -7091 37 -7075 71
rect -6987 37 -6971 71
rect -6913 37 -6897 71
rect -6809 37 -6793 71
rect -6735 37 -6719 71
rect -6631 37 -6615 71
rect -6557 37 -6541 71
rect -6453 37 -6437 71
rect -6379 37 -6363 71
rect -6275 37 -6259 71
rect -6201 37 -6185 71
rect -6097 37 -6081 71
rect -6023 37 -6007 71
rect -5919 37 -5903 71
rect -5845 37 -5829 71
rect -5741 37 -5725 71
rect -5667 37 -5651 71
rect -5563 37 -5547 71
rect -5489 37 -5473 71
rect -5385 37 -5369 71
rect -5311 37 -5295 71
rect -5207 37 -5191 71
rect -5133 37 -5117 71
rect -5029 37 -5013 71
rect -4955 37 -4939 71
rect -4851 37 -4835 71
rect -4777 37 -4761 71
rect -4673 37 -4657 71
rect -4599 37 -4583 71
rect -4495 37 -4479 71
rect -4421 37 -4405 71
rect -4317 37 -4301 71
rect -4243 37 -4227 71
rect -4139 37 -4123 71
rect -4065 37 -4049 71
rect -3961 37 -3945 71
rect -3887 37 -3871 71
rect -3783 37 -3767 71
rect -3709 37 -3693 71
rect -3605 37 -3589 71
rect -3531 37 -3515 71
rect -3427 37 -3411 71
rect -3353 37 -3337 71
rect -3249 37 -3233 71
rect -3175 37 -3159 71
rect -3071 37 -3055 71
rect -2997 37 -2981 71
rect -2893 37 -2877 71
rect -2819 37 -2803 71
rect -2715 37 -2699 71
rect -2641 37 -2625 71
rect -2537 37 -2521 71
rect -2463 37 -2447 71
rect -2359 37 -2343 71
rect -2285 37 -2269 71
rect -2181 37 -2165 71
rect -2107 37 -2091 71
rect -2003 37 -1987 71
rect -1929 37 -1913 71
rect -1825 37 -1809 71
rect -1751 37 -1735 71
rect -1647 37 -1631 71
rect -1573 37 -1557 71
rect -1469 37 -1453 71
rect -1395 37 -1379 71
rect -1291 37 -1275 71
rect -1217 37 -1201 71
rect -1113 37 -1097 71
rect -1039 37 -1023 71
rect -935 37 -919 71
rect -861 37 -845 71
rect -757 37 -741 71
rect -683 37 -667 71
rect -579 37 -563 71
rect -505 37 -489 71
rect -401 37 -385 71
rect -327 37 -311 71
rect -223 37 -207 71
rect -149 37 -133 71
rect -45 37 -29 71
rect 29 37 45 71
rect 133 37 149 71
rect 207 37 223 71
rect 311 37 327 71
rect 385 37 401 71
rect 489 37 505 71
rect 563 37 579 71
rect 667 37 683 71
rect 741 37 757 71
rect 845 37 861 71
rect 919 37 935 71
rect 1023 37 1039 71
rect 1097 37 1113 71
rect 1201 37 1217 71
rect 1275 37 1291 71
rect 1379 37 1395 71
rect 1453 37 1469 71
rect 1557 37 1573 71
rect 1631 37 1647 71
rect 1735 37 1751 71
rect 1809 37 1825 71
rect 1913 37 1929 71
rect 1987 37 2003 71
rect 2091 37 2107 71
rect 2165 37 2181 71
rect 2269 37 2285 71
rect 2343 37 2359 71
rect 2447 37 2463 71
rect 2521 37 2537 71
rect 2625 37 2641 71
rect 2699 37 2715 71
rect 2803 37 2819 71
rect 2877 37 2893 71
rect 2981 37 2997 71
rect 3055 37 3071 71
rect 3159 37 3175 71
rect 3233 37 3249 71
rect 3337 37 3353 71
rect 3411 37 3427 71
rect 3515 37 3531 71
rect 3589 37 3605 71
rect 3693 37 3709 71
rect 3767 37 3783 71
rect 3871 37 3887 71
rect 3945 37 3961 71
rect 4049 37 4065 71
rect 4123 37 4139 71
rect 4227 37 4243 71
rect 4301 37 4317 71
rect 4405 37 4421 71
rect 4479 37 4495 71
rect 4583 37 4599 71
rect 4657 37 4673 71
rect 4761 37 4777 71
rect 4835 37 4851 71
rect 4939 37 4955 71
rect 5013 37 5029 71
rect 5117 37 5133 71
rect 5191 37 5207 71
rect 5295 37 5311 71
rect 5369 37 5385 71
rect 5473 37 5489 71
rect 5547 37 5563 71
rect 5651 37 5667 71
rect 5725 37 5741 71
rect 5829 37 5845 71
rect 5903 37 5919 71
rect 6007 37 6023 71
rect 6081 37 6097 71
rect 6185 37 6201 71
rect 6259 37 6275 71
rect 6363 37 6379 71
rect 6437 37 6453 71
rect 6541 37 6557 71
rect 6615 37 6631 71
rect 6719 37 6735 71
rect 6793 37 6809 71
rect 6897 37 6913 71
rect 6971 37 6987 71
rect 7075 37 7091 71
rect 7149 37 7165 71
rect 7253 37 7269 71
rect 7327 37 7343 71
rect 7431 37 7447 71
rect 7505 37 7521 71
rect 7609 37 7625 71
rect 7683 37 7699 71
rect 7787 37 7803 71
rect 7861 37 7877 71
rect 7965 37 7981 71
rect 8039 37 8055 71
rect 8143 37 8159 71
rect 8217 37 8233 71
rect 8321 37 8337 71
rect 8395 37 8411 71
rect 8499 37 8515 71
rect 8573 37 8589 71
rect 8677 37 8693 71
rect 8751 37 8767 71
rect 8855 37 8871 71
rect -8871 -71 -8855 -37
rect -8767 -71 -8751 -37
rect -8693 -71 -8677 -37
rect -8589 -71 -8573 -37
rect -8515 -71 -8499 -37
rect -8411 -71 -8395 -37
rect -8337 -71 -8321 -37
rect -8233 -71 -8217 -37
rect -8159 -71 -8143 -37
rect -8055 -71 -8039 -37
rect -7981 -71 -7965 -37
rect -7877 -71 -7861 -37
rect -7803 -71 -7787 -37
rect -7699 -71 -7683 -37
rect -7625 -71 -7609 -37
rect -7521 -71 -7505 -37
rect -7447 -71 -7431 -37
rect -7343 -71 -7327 -37
rect -7269 -71 -7253 -37
rect -7165 -71 -7149 -37
rect -7091 -71 -7075 -37
rect -6987 -71 -6971 -37
rect -6913 -71 -6897 -37
rect -6809 -71 -6793 -37
rect -6735 -71 -6719 -37
rect -6631 -71 -6615 -37
rect -6557 -71 -6541 -37
rect -6453 -71 -6437 -37
rect -6379 -71 -6363 -37
rect -6275 -71 -6259 -37
rect -6201 -71 -6185 -37
rect -6097 -71 -6081 -37
rect -6023 -71 -6007 -37
rect -5919 -71 -5903 -37
rect -5845 -71 -5829 -37
rect -5741 -71 -5725 -37
rect -5667 -71 -5651 -37
rect -5563 -71 -5547 -37
rect -5489 -71 -5473 -37
rect -5385 -71 -5369 -37
rect -5311 -71 -5295 -37
rect -5207 -71 -5191 -37
rect -5133 -71 -5117 -37
rect -5029 -71 -5013 -37
rect -4955 -71 -4939 -37
rect -4851 -71 -4835 -37
rect -4777 -71 -4761 -37
rect -4673 -71 -4657 -37
rect -4599 -71 -4583 -37
rect -4495 -71 -4479 -37
rect -4421 -71 -4405 -37
rect -4317 -71 -4301 -37
rect -4243 -71 -4227 -37
rect -4139 -71 -4123 -37
rect -4065 -71 -4049 -37
rect -3961 -71 -3945 -37
rect -3887 -71 -3871 -37
rect -3783 -71 -3767 -37
rect -3709 -71 -3693 -37
rect -3605 -71 -3589 -37
rect -3531 -71 -3515 -37
rect -3427 -71 -3411 -37
rect -3353 -71 -3337 -37
rect -3249 -71 -3233 -37
rect -3175 -71 -3159 -37
rect -3071 -71 -3055 -37
rect -2997 -71 -2981 -37
rect -2893 -71 -2877 -37
rect -2819 -71 -2803 -37
rect -2715 -71 -2699 -37
rect -2641 -71 -2625 -37
rect -2537 -71 -2521 -37
rect -2463 -71 -2447 -37
rect -2359 -71 -2343 -37
rect -2285 -71 -2269 -37
rect -2181 -71 -2165 -37
rect -2107 -71 -2091 -37
rect -2003 -71 -1987 -37
rect -1929 -71 -1913 -37
rect -1825 -71 -1809 -37
rect -1751 -71 -1735 -37
rect -1647 -71 -1631 -37
rect -1573 -71 -1557 -37
rect -1469 -71 -1453 -37
rect -1395 -71 -1379 -37
rect -1291 -71 -1275 -37
rect -1217 -71 -1201 -37
rect -1113 -71 -1097 -37
rect -1039 -71 -1023 -37
rect -935 -71 -919 -37
rect -861 -71 -845 -37
rect -757 -71 -741 -37
rect -683 -71 -667 -37
rect -579 -71 -563 -37
rect -505 -71 -489 -37
rect -401 -71 -385 -37
rect -327 -71 -311 -37
rect -223 -71 -207 -37
rect -149 -71 -133 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 133 -71 149 -37
rect 207 -71 223 -37
rect 311 -71 327 -37
rect 385 -71 401 -37
rect 489 -71 505 -37
rect 563 -71 579 -37
rect 667 -71 683 -37
rect 741 -71 757 -37
rect 845 -71 861 -37
rect 919 -71 935 -37
rect 1023 -71 1039 -37
rect 1097 -71 1113 -37
rect 1201 -71 1217 -37
rect 1275 -71 1291 -37
rect 1379 -71 1395 -37
rect 1453 -71 1469 -37
rect 1557 -71 1573 -37
rect 1631 -71 1647 -37
rect 1735 -71 1751 -37
rect 1809 -71 1825 -37
rect 1913 -71 1929 -37
rect 1987 -71 2003 -37
rect 2091 -71 2107 -37
rect 2165 -71 2181 -37
rect 2269 -71 2285 -37
rect 2343 -71 2359 -37
rect 2447 -71 2463 -37
rect 2521 -71 2537 -37
rect 2625 -71 2641 -37
rect 2699 -71 2715 -37
rect 2803 -71 2819 -37
rect 2877 -71 2893 -37
rect 2981 -71 2997 -37
rect 3055 -71 3071 -37
rect 3159 -71 3175 -37
rect 3233 -71 3249 -37
rect 3337 -71 3353 -37
rect 3411 -71 3427 -37
rect 3515 -71 3531 -37
rect 3589 -71 3605 -37
rect 3693 -71 3709 -37
rect 3767 -71 3783 -37
rect 3871 -71 3887 -37
rect 3945 -71 3961 -37
rect 4049 -71 4065 -37
rect 4123 -71 4139 -37
rect 4227 -71 4243 -37
rect 4301 -71 4317 -37
rect 4405 -71 4421 -37
rect 4479 -71 4495 -37
rect 4583 -71 4599 -37
rect 4657 -71 4673 -37
rect 4761 -71 4777 -37
rect 4835 -71 4851 -37
rect 4939 -71 4955 -37
rect 5013 -71 5029 -37
rect 5117 -71 5133 -37
rect 5191 -71 5207 -37
rect 5295 -71 5311 -37
rect 5369 -71 5385 -37
rect 5473 -71 5489 -37
rect 5547 -71 5563 -37
rect 5651 -71 5667 -37
rect 5725 -71 5741 -37
rect 5829 -71 5845 -37
rect 5903 -71 5919 -37
rect 6007 -71 6023 -37
rect 6081 -71 6097 -37
rect 6185 -71 6201 -37
rect 6259 -71 6275 -37
rect 6363 -71 6379 -37
rect 6437 -71 6453 -37
rect 6541 -71 6557 -37
rect 6615 -71 6631 -37
rect 6719 -71 6735 -37
rect 6793 -71 6809 -37
rect 6897 -71 6913 -37
rect 6971 -71 6987 -37
rect 7075 -71 7091 -37
rect 7149 -71 7165 -37
rect 7253 -71 7269 -37
rect 7327 -71 7343 -37
rect 7431 -71 7447 -37
rect 7505 -71 7521 -37
rect 7609 -71 7625 -37
rect 7683 -71 7699 -37
rect 7787 -71 7803 -37
rect 7861 -71 7877 -37
rect 7965 -71 7981 -37
rect 8039 -71 8055 -37
rect 8143 -71 8159 -37
rect 8217 -71 8233 -37
rect 8321 -71 8337 -37
rect 8395 -71 8411 -37
rect 8499 -71 8515 -37
rect 8573 -71 8589 -37
rect 8677 -71 8693 -37
rect 8751 -71 8767 -37
rect 8855 -71 8871 -37
rect -8917 -130 -8883 -114
rect -8917 -2522 -8883 -2506
rect -8739 -130 -8705 -114
rect -8739 -2522 -8705 -2506
rect -8561 -130 -8527 -114
rect -8561 -2522 -8527 -2506
rect -8383 -130 -8349 -114
rect -8383 -2522 -8349 -2506
rect -8205 -130 -8171 -114
rect -8205 -2522 -8171 -2506
rect -8027 -130 -7993 -114
rect -8027 -2522 -7993 -2506
rect -7849 -130 -7815 -114
rect -7849 -2522 -7815 -2506
rect -7671 -130 -7637 -114
rect -7671 -2522 -7637 -2506
rect -7493 -130 -7459 -114
rect -7493 -2522 -7459 -2506
rect -7315 -130 -7281 -114
rect -7315 -2522 -7281 -2506
rect -7137 -130 -7103 -114
rect -7137 -2522 -7103 -2506
rect -6959 -130 -6925 -114
rect -6959 -2522 -6925 -2506
rect -6781 -130 -6747 -114
rect -6781 -2522 -6747 -2506
rect -6603 -130 -6569 -114
rect -6603 -2522 -6569 -2506
rect -6425 -130 -6391 -114
rect -6425 -2522 -6391 -2506
rect -6247 -130 -6213 -114
rect -6247 -2522 -6213 -2506
rect -6069 -130 -6035 -114
rect -6069 -2522 -6035 -2506
rect -5891 -130 -5857 -114
rect -5891 -2522 -5857 -2506
rect -5713 -130 -5679 -114
rect -5713 -2522 -5679 -2506
rect -5535 -130 -5501 -114
rect -5535 -2522 -5501 -2506
rect -5357 -130 -5323 -114
rect -5357 -2522 -5323 -2506
rect -5179 -130 -5145 -114
rect -5179 -2522 -5145 -2506
rect -5001 -130 -4967 -114
rect -5001 -2522 -4967 -2506
rect -4823 -130 -4789 -114
rect -4823 -2522 -4789 -2506
rect -4645 -130 -4611 -114
rect -4645 -2522 -4611 -2506
rect -4467 -130 -4433 -114
rect -4467 -2522 -4433 -2506
rect -4289 -130 -4255 -114
rect -4289 -2522 -4255 -2506
rect -4111 -130 -4077 -114
rect -4111 -2522 -4077 -2506
rect -3933 -130 -3899 -114
rect -3933 -2522 -3899 -2506
rect -3755 -130 -3721 -114
rect -3755 -2522 -3721 -2506
rect -3577 -130 -3543 -114
rect -3577 -2522 -3543 -2506
rect -3399 -130 -3365 -114
rect -3399 -2522 -3365 -2506
rect -3221 -130 -3187 -114
rect -3221 -2522 -3187 -2506
rect -3043 -130 -3009 -114
rect -3043 -2522 -3009 -2506
rect -2865 -130 -2831 -114
rect -2865 -2522 -2831 -2506
rect -2687 -130 -2653 -114
rect -2687 -2522 -2653 -2506
rect -2509 -130 -2475 -114
rect -2509 -2522 -2475 -2506
rect -2331 -130 -2297 -114
rect -2331 -2522 -2297 -2506
rect -2153 -130 -2119 -114
rect -2153 -2522 -2119 -2506
rect -1975 -130 -1941 -114
rect -1975 -2522 -1941 -2506
rect -1797 -130 -1763 -114
rect -1797 -2522 -1763 -2506
rect -1619 -130 -1585 -114
rect -1619 -2522 -1585 -2506
rect -1441 -130 -1407 -114
rect -1441 -2522 -1407 -2506
rect -1263 -130 -1229 -114
rect -1263 -2522 -1229 -2506
rect -1085 -130 -1051 -114
rect -1085 -2522 -1051 -2506
rect -907 -130 -873 -114
rect -907 -2522 -873 -2506
rect -729 -130 -695 -114
rect -729 -2522 -695 -2506
rect -551 -130 -517 -114
rect -551 -2522 -517 -2506
rect -373 -130 -339 -114
rect -373 -2522 -339 -2506
rect -195 -130 -161 -114
rect -195 -2522 -161 -2506
rect -17 -130 17 -114
rect -17 -2522 17 -2506
rect 161 -130 195 -114
rect 161 -2522 195 -2506
rect 339 -130 373 -114
rect 339 -2522 373 -2506
rect 517 -130 551 -114
rect 517 -2522 551 -2506
rect 695 -130 729 -114
rect 695 -2522 729 -2506
rect 873 -130 907 -114
rect 873 -2522 907 -2506
rect 1051 -130 1085 -114
rect 1051 -2522 1085 -2506
rect 1229 -130 1263 -114
rect 1229 -2522 1263 -2506
rect 1407 -130 1441 -114
rect 1407 -2522 1441 -2506
rect 1585 -130 1619 -114
rect 1585 -2522 1619 -2506
rect 1763 -130 1797 -114
rect 1763 -2522 1797 -2506
rect 1941 -130 1975 -114
rect 1941 -2522 1975 -2506
rect 2119 -130 2153 -114
rect 2119 -2522 2153 -2506
rect 2297 -130 2331 -114
rect 2297 -2522 2331 -2506
rect 2475 -130 2509 -114
rect 2475 -2522 2509 -2506
rect 2653 -130 2687 -114
rect 2653 -2522 2687 -2506
rect 2831 -130 2865 -114
rect 2831 -2522 2865 -2506
rect 3009 -130 3043 -114
rect 3009 -2522 3043 -2506
rect 3187 -130 3221 -114
rect 3187 -2522 3221 -2506
rect 3365 -130 3399 -114
rect 3365 -2522 3399 -2506
rect 3543 -130 3577 -114
rect 3543 -2522 3577 -2506
rect 3721 -130 3755 -114
rect 3721 -2522 3755 -2506
rect 3899 -130 3933 -114
rect 3899 -2522 3933 -2506
rect 4077 -130 4111 -114
rect 4077 -2522 4111 -2506
rect 4255 -130 4289 -114
rect 4255 -2522 4289 -2506
rect 4433 -130 4467 -114
rect 4433 -2522 4467 -2506
rect 4611 -130 4645 -114
rect 4611 -2522 4645 -2506
rect 4789 -130 4823 -114
rect 4789 -2522 4823 -2506
rect 4967 -130 5001 -114
rect 4967 -2522 5001 -2506
rect 5145 -130 5179 -114
rect 5145 -2522 5179 -2506
rect 5323 -130 5357 -114
rect 5323 -2522 5357 -2506
rect 5501 -130 5535 -114
rect 5501 -2522 5535 -2506
rect 5679 -130 5713 -114
rect 5679 -2522 5713 -2506
rect 5857 -130 5891 -114
rect 5857 -2522 5891 -2506
rect 6035 -130 6069 -114
rect 6035 -2522 6069 -2506
rect 6213 -130 6247 -114
rect 6213 -2522 6247 -2506
rect 6391 -130 6425 -114
rect 6391 -2522 6425 -2506
rect 6569 -130 6603 -114
rect 6569 -2522 6603 -2506
rect 6747 -130 6781 -114
rect 6747 -2522 6781 -2506
rect 6925 -130 6959 -114
rect 6925 -2522 6959 -2506
rect 7103 -130 7137 -114
rect 7103 -2522 7137 -2506
rect 7281 -130 7315 -114
rect 7281 -2522 7315 -2506
rect 7459 -130 7493 -114
rect 7459 -2522 7493 -2506
rect 7637 -130 7671 -114
rect 7637 -2522 7671 -2506
rect 7815 -130 7849 -114
rect 7815 -2522 7849 -2506
rect 7993 -130 8027 -114
rect 7993 -2522 8027 -2506
rect 8171 -130 8205 -114
rect 8171 -2522 8205 -2506
rect 8349 -130 8383 -114
rect 8349 -2522 8383 -2506
rect 8527 -130 8561 -114
rect 8527 -2522 8561 -2506
rect 8705 -130 8739 -114
rect 8705 -2522 8739 -2506
rect 8883 -130 8917 -114
rect 8883 -2522 8917 -2506
rect -8871 -2599 -8855 -2565
rect -8767 -2599 -8751 -2565
rect -8693 -2599 -8677 -2565
rect -8589 -2599 -8573 -2565
rect -8515 -2599 -8499 -2565
rect -8411 -2599 -8395 -2565
rect -8337 -2599 -8321 -2565
rect -8233 -2599 -8217 -2565
rect -8159 -2599 -8143 -2565
rect -8055 -2599 -8039 -2565
rect -7981 -2599 -7965 -2565
rect -7877 -2599 -7861 -2565
rect -7803 -2599 -7787 -2565
rect -7699 -2599 -7683 -2565
rect -7625 -2599 -7609 -2565
rect -7521 -2599 -7505 -2565
rect -7447 -2599 -7431 -2565
rect -7343 -2599 -7327 -2565
rect -7269 -2599 -7253 -2565
rect -7165 -2599 -7149 -2565
rect -7091 -2599 -7075 -2565
rect -6987 -2599 -6971 -2565
rect -6913 -2599 -6897 -2565
rect -6809 -2599 -6793 -2565
rect -6735 -2599 -6719 -2565
rect -6631 -2599 -6615 -2565
rect -6557 -2599 -6541 -2565
rect -6453 -2599 -6437 -2565
rect -6379 -2599 -6363 -2565
rect -6275 -2599 -6259 -2565
rect -6201 -2599 -6185 -2565
rect -6097 -2599 -6081 -2565
rect -6023 -2599 -6007 -2565
rect -5919 -2599 -5903 -2565
rect -5845 -2599 -5829 -2565
rect -5741 -2599 -5725 -2565
rect -5667 -2599 -5651 -2565
rect -5563 -2599 -5547 -2565
rect -5489 -2599 -5473 -2565
rect -5385 -2599 -5369 -2565
rect -5311 -2599 -5295 -2565
rect -5207 -2599 -5191 -2565
rect -5133 -2599 -5117 -2565
rect -5029 -2599 -5013 -2565
rect -4955 -2599 -4939 -2565
rect -4851 -2599 -4835 -2565
rect -4777 -2599 -4761 -2565
rect -4673 -2599 -4657 -2565
rect -4599 -2599 -4583 -2565
rect -4495 -2599 -4479 -2565
rect -4421 -2599 -4405 -2565
rect -4317 -2599 -4301 -2565
rect -4243 -2599 -4227 -2565
rect -4139 -2599 -4123 -2565
rect -4065 -2599 -4049 -2565
rect -3961 -2599 -3945 -2565
rect -3887 -2599 -3871 -2565
rect -3783 -2599 -3767 -2565
rect -3709 -2599 -3693 -2565
rect -3605 -2599 -3589 -2565
rect -3531 -2599 -3515 -2565
rect -3427 -2599 -3411 -2565
rect -3353 -2599 -3337 -2565
rect -3249 -2599 -3233 -2565
rect -3175 -2599 -3159 -2565
rect -3071 -2599 -3055 -2565
rect -2997 -2599 -2981 -2565
rect -2893 -2599 -2877 -2565
rect -2819 -2599 -2803 -2565
rect -2715 -2599 -2699 -2565
rect -2641 -2599 -2625 -2565
rect -2537 -2599 -2521 -2565
rect -2463 -2599 -2447 -2565
rect -2359 -2599 -2343 -2565
rect -2285 -2599 -2269 -2565
rect -2181 -2599 -2165 -2565
rect -2107 -2599 -2091 -2565
rect -2003 -2599 -1987 -2565
rect -1929 -2599 -1913 -2565
rect -1825 -2599 -1809 -2565
rect -1751 -2599 -1735 -2565
rect -1647 -2599 -1631 -2565
rect -1573 -2599 -1557 -2565
rect -1469 -2599 -1453 -2565
rect -1395 -2599 -1379 -2565
rect -1291 -2599 -1275 -2565
rect -1217 -2599 -1201 -2565
rect -1113 -2599 -1097 -2565
rect -1039 -2599 -1023 -2565
rect -935 -2599 -919 -2565
rect -861 -2599 -845 -2565
rect -757 -2599 -741 -2565
rect -683 -2599 -667 -2565
rect -579 -2599 -563 -2565
rect -505 -2599 -489 -2565
rect -401 -2599 -385 -2565
rect -327 -2599 -311 -2565
rect -223 -2599 -207 -2565
rect -149 -2599 -133 -2565
rect -45 -2599 -29 -2565
rect 29 -2599 45 -2565
rect 133 -2599 149 -2565
rect 207 -2599 223 -2565
rect 311 -2599 327 -2565
rect 385 -2599 401 -2565
rect 489 -2599 505 -2565
rect 563 -2599 579 -2565
rect 667 -2599 683 -2565
rect 741 -2599 757 -2565
rect 845 -2599 861 -2565
rect 919 -2599 935 -2565
rect 1023 -2599 1039 -2565
rect 1097 -2599 1113 -2565
rect 1201 -2599 1217 -2565
rect 1275 -2599 1291 -2565
rect 1379 -2599 1395 -2565
rect 1453 -2599 1469 -2565
rect 1557 -2599 1573 -2565
rect 1631 -2599 1647 -2565
rect 1735 -2599 1751 -2565
rect 1809 -2599 1825 -2565
rect 1913 -2599 1929 -2565
rect 1987 -2599 2003 -2565
rect 2091 -2599 2107 -2565
rect 2165 -2599 2181 -2565
rect 2269 -2599 2285 -2565
rect 2343 -2599 2359 -2565
rect 2447 -2599 2463 -2565
rect 2521 -2599 2537 -2565
rect 2625 -2599 2641 -2565
rect 2699 -2599 2715 -2565
rect 2803 -2599 2819 -2565
rect 2877 -2599 2893 -2565
rect 2981 -2599 2997 -2565
rect 3055 -2599 3071 -2565
rect 3159 -2599 3175 -2565
rect 3233 -2599 3249 -2565
rect 3337 -2599 3353 -2565
rect 3411 -2599 3427 -2565
rect 3515 -2599 3531 -2565
rect 3589 -2599 3605 -2565
rect 3693 -2599 3709 -2565
rect 3767 -2599 3783 -2565
rect 3871 -2599 3887 -2565
rect 3945 -2599 3961 -2565
rect 4049 -2599 4065 -2565
rect 4123 -2599 4139 -2565
rect 4227 -2599 4243 -2565
rect 4301 -2599 4317 -2565
rect 4405 -2599 4421 -2565
rect 4479 -2599 4495 -2565
rect 4583 -2599 4599 -2565
rect 4657 -2599 4673 -2565
rect 4761 -2599 4777 -2565
rect 4835 -2599 4851 -2565
rect 4939 -2599 4955 -2565
rect 5013 -2599 5029 -2565
rect 5117 -2599 5133 -2565
rect 5191 -2599 5207 -2565
rect 5295 -2599 5311 -2565
rect 5369 -2599 5385 -2565
rect 5473 -2599 5489 -2565
rect 5547 -2599 5563 -2565
rect 5651 -2599 5667 -2565
rect 5725 -2599 5741 -2565
rect 5829 -2599 5845 -2565
rect 5903 -2599 5919 -2565
rect 6007 -2599 6023 -2565
rect 6081 -2599 6097 -2565
rect 6185 -2599 6201 -2565
rect 6259 -2599 6275 -2565
rect 6363 -2599 6379 -2565
rect 6437 -2599 6453 -2565
rect 6541 -2599 6557 -2565
rect 6615 -2599 6631 -2565
rect 6719 -2599 6735 -2565
rect 6793 -2599 6809 -2565
rect 6897 -2599 6913 -2565
rect 6971 -2599 6987 -2565
rect 7075 -2599 7091 -2565
rect 7149 -2599 7165 -2565
rect 7253 -2599 7269 -2565
rect 7327 -2599 7343 -2565
rect 7431 -2599 7447 -2565
rect 7505 -2599 7521 -2565
rect 7609 -2599 7625 -2565
rect 7683 -2599 7699 -2565
rect 7787 -2599 7803 -2565
rect 7861 -2599 7877 -2565
rect 7965 -2599 7981 -2565
rect 8039 -2599 8055 -2565
rect 8143 -2599 8159 -2565
rect 8217 -2599 8233 -2565
rect 8321 -2599 8337 -2565
rect 8395 -2599 8411 -2565
rect 8499 -2599 8515 -2565
rect 8573 -2599 8589 -2565
rect 8677 -2599 8693 -2565
rect 8751 -2599 8767 -2565
rect 8855 -2599 8871 -2565
rect -9031 -2667 -8997 -2605
rect 8997 -2667 9031 -2605
rect -9031 -2701 -8935 -2667
rect 8935 -2701 9031 -2667
<< viali >>
rect -8855 2565 -8767 2599
rect -8677 2565 -8589 2599
rect -8499 2565 -8411 2599
rect -8321 2565 -8233 2599
rect -8143 2565 -8055 2599
rect -7965 2565 -7877 2599
rect -7787 2565 -7699 2599
rect -7609 2565 -7521 2599
rect -7431 2565 -7343 2599
rect -7253 2565 -7165 2599
rect -7075 2565 -6987 2599
rect -6897 2565 -6809 2599
rect -6719 2565 -6631 2599
rect -6541 2565 -6453 2599
rect -6363 2565 -6275 2599
rect -6185 2565 -6097 2599
rect -6007 2565 -5919 2599
rect -5829 2565 -5741 2599
rect -5651 2565 -5563 2599
rect -5473 2565 -5385 2599
rect -5295 2565 -5207 2599
rect -5117 2565 -5029 2599
rect -4939 2565 -4851 2599
rect -4761 2565 -4673 2599
rect -4583 2565 -4495 2599
rect -4405 2565 -4317 2599
rect -4227 2565 -4139 2599
rect -4049 2565 -3961 2599
rect -3871 2565 -3783 2599
rect -3693 2565 -3605 2599
rect -3515 2565 -3427 2599
rect -3337 2565 -3249 2599
rect -3159 2565 -3071 2599
rect -2981 2565 -2893 2599
rect -2803 2565 -2715 2599
rect -2625 2565 -2537 2599
rect -2447 2565 -2359 2599
rect -2269 2565 -2181 2599
rect -2091 2565 -2003 2599
rect -1913 2565 -1825 2599
rect -1735 2565 -1647 2599
rect -1557 2565 -1469 2599
rect -1379 2565 -1291 2599
rect -1201 2565 -1113 2599
rect -1023 2565 -935 2599
rect -845 2565 -757 2599
rect -667 2565 -579 2599
rect -489 2565 -401 2599
rect -311 2565 -223 2599
rect -133 2565 -45 2599
rect 45 2565 133 2599
rect 223 2565 311 2599
rect 401 2565 489 2599
rect 579 2565 667 2599
rect 757 2565 845 2599
rect 935 2565 1023 2599
rect 1113 2565 1201 2599
rect 1291 2565 1379 2599
rect 1469 2565 1557 2599
rect 1647 2565 1735 2599
rect 1825 2565 1913 2599
rect 2003 2565 2091 2599
rect 2181 2565 2269 2599
rect 2359 2565 2447 2599
rect 2537 2565 2625 2599
rect 2715 2565 2803 2599
rect 2893 2565 2981 2599
rect 3071 2565 3159 2599
rect 3249 2565 3337 2599
rect 3427 2565 3515 2599
rect 3605 2565 3693 2599
rect 3783 2565 3871 2599
rect 3961 2565 4049 2599
rect 4139 2565 4227 2599
rect 4317 2565 4405 2599
rect 4495 2565 4583 2599
rect 4673 2565 4761 2599
rect 4851 2565 4939 2599
rect 5029 2565 5117 2599
rect 5207 2565 5295 2599
rect 5385 2565 5473 2599
rect 5563 2565 5651 2599
rect 5741 2565 5829 2599
rect 5919 2565 6007 2599
rect 6097 2565 6185 2599
rect 6275 2565 6363 2599
rect 6453 2565 6541 2599
rect 6631 2565 6719 2599
rect 6809 2565 6897 2599
rect 6987 2565 7075 2599
rect 7165 2565 7253 2599
rect 7343 2565 7431 2599
rect 7521 2565 7609 2599
rect 7699 2565 7787 2599
rect 7877 2565 7965 2599
rect 8055 2565 8143 2599
rect 8233 2565 8321 2599
rect 8411 2565 8499 2599
rect 8589 2565 8677 2599
rect 8767 2565 8855 2599
rect -8917 130 -8883 2506
rect -8739 130 -8705 2506
rect -8561 130 -8527 2506
rect -8383 130 -8349 2506
rect -8205 130 -8171 2506
rect -8027 130 -7993 2506
rect -7849 130 -7815 2506
rect -7671 130 -7637 2506
rect -7493 130 -7459 2506
rect -7315 130 -7281 2506
rect -7137 130 -7103 2506
rect -6959 130 -6925 2506
rect -6781 130 -6747 2506
rect -6603 130 -6569 2506
rect -6425 130 -6391 2506
rect -6247 130 -6213 2506
rect -6069 130 -6035 2506
rect -5891 130 -5857 2506
rect -5713 130 -5679 2506
rect -5535 130 -5501 2506
rect -5357 130 -5323 2506
rect -5179 130 -5145 2506
rect -5001 130 -4967 2506
rect -4823 130 -4789 2506
rect -4645 130 -4611 2506
rect -4467 130 -4433 2506
rect -4289 130 -4255 2506
rect -4111 130 -4077 2506
rect -3933 130 -3899 2506
rect -3755 130 -3721 2506
rect -3577 130 -3543 2506
rect -3399 130 -3365 2506
rect -3221 130 -3187 2506
rect -3043 130 -3009 2506
rect -2865 130 -2831 2506
rect -2687 130 -2653 2506
rect -2509 130 -2475 2506
rect -2331 130 -2297 2506
rect -2153 130 -2119 2506
rect -1975 130 -1941 2506
rect -1797 130 -1763 2506
rect -1619 130 -1585 2506
rect -1441 130 -1407 2506
rect -1263 130 -1229 2506
rect -1085 130 -1051 2506
rect -907 130 -873 2506
rect -729 130 -695 2506
rect -551 130 -517 2506
rect -373 130 -339 2506
rect -195 130 -161 2506
rect -17 130 17 2506
rect 161 130 195 2506
rect 339 130 373 2506
rect 517 130 551 2506
rect 695 130 729 2506
rect 873 130 907 2506
rect 1051 130 1085 2506
rect 1229 130 1263 2506
rect 1407 130 1441 2506
rect 1585 130 1619 2506
rect 1763 130 1797 2506
rect 1941 130 1975 2506
rect 2119 130 2153 2506
rect 2297 130 2331 2506
rect 2475 130 2509 2506
rect 2653 130 2687 2506
rect 2831 130 2865 2506
rect 3009 130 3043 2506
rect 3187 130 3221 2506
rect 3365 130 3399 2506
rect 3543 130 3577 2506
rect 3721 130 3755 2506
rect 3899 130 3933 2506
rect 4077 130 4111 2506
rect 4255 130 4289 2506
rect 4433 130 4467 2506
rect 4611 130 4645 2506
rect 4789 130 4823 2506
rect 4967 130 5001 2506
rect 5145 130 5179 2506
rect 5323 130 5357 2506
rect 5501 130 5535 2506
rect 5679 130 5713 2506
rect 5857 130 5891 2506
rect 6035 130 6069 2506
rect 6213 130 6247 2506
rect 6391 130 6425 2506
rect 6569 130 6603 2506
rect 6747 130 6781 2506
rect 6925 130 6959 2506
rect 7103 130 7137 2506
rect 7281 130 7315 2506
rect 7459 130 7493 2506
rect 7637 130 7671 2506
rect 7815 130 7849 2506
rect 7993 130 8027 2506
rect 8171 130 8205 2506
rect 8349 130 8383 2506
rect 8527 130 8561 2506
rect 8705 130 8739 2506
rect 8883 130 8917 2506
rect -8855 37 -8767 71
rect -8677 37 -8589 71
rect -8499 37 -8411 71
rect -8321 37 -8233 71
rect -8143 37 -8055 71
rect -7965 37 -7877 71
rect -7787 37 -7699 71
rect -7609 37 -7521 71
rect -7431 37 -7343 71
rect -7253 37 -7165 71
rect -7075 37 -6987 71
rect -6897 37 -6809 71
rect -6719 37 -6631 71
rect -6541 37 -6453 71
rect -6363 37 -6275 71
rect -6185 37 -6097 71
rect -6007 37 -5919 71
rect -5829 37 -5741 71
rect -5651 37 -5563 71
rect -5473 37 -5385 71
rect -5295 37 -5207 71
rect -5117 37 -5029 71
rect -4939 37 -4851 71
rect -4761 37 -4673 71
rect -4583 37 -4495 71
rect -4405 37 -4317 71
rect -4227 37 -4139 71
rect -4049 37 -3961 71
rect -3871 37 -3783 71
rect -3693 37 -3605 71
rect -3515 37 -3427 71
rect -3337 37 -3249 71
rect -3159 37 -3071 71
rect -2981 37 -2893 71
rect -2803 37 -2715 71
rect -2625 37 -2537 71
rect -2447 37 -2359 71
rect -2269 37 -2181 71
rect -2091 37 -2003 71
rect -1913 37 -1825 71
rect -1735 37 -1647 71
rect -1557 37 -1469 71
rect -1379 37 -1291 71
rect -1201 37 -1113 71
rect -1023 37 -935 71
rect -845 37 -757 71
rect -667 37 -579 71
rect -489 37 -401 71
rect -311 37 -223 71
rect -133 37 -45 71
rect 45 37 133 71
rect 223 37 311 71
rect 401 37 489 71
rect 579 37 667 71
rect 757 37 845 71
rect 935 37 1023 71
rect 1113 37 1201 71
rect 1291 37 1379 71
rect 1469 37 1557 71
rect 1647 37 1735 71
rect 1825 37 1913 71
rect 2003 37 2091 71
rect 2181 37 2269 71
rect 2359 37 2447 71
rect 2537 37 2625 71
rect 2715 37 2803 71
rect 2893 37 2981 71
rect 3071 37 3159 71
rect 3249 37 3337 71
rect 3427 37 3515 71
rect 3605 37 3693 71
rect 3783 37 3871 71
rect 3961 37 4049 71
rect 4139 37 4227 71
rect 4317 37 4405 71
rect 4495 37 4583 71
rect 4673 37 4761 71
rect 4851 37 4939 71
rect 5029 37 5117 71
rect 5207 37 5295 71
rect 5385 37 5473 71
rect 5563 37 5651 71
rect 5741 37 5829 71
rect 5919 37 6007 71
rect 6097 37 6185 71
rect 6275 37 6363 71
rect 6453 37 6541 71
rect 6631 37 6719 71
rect 6809 37 6897 71
rect 6987 37 7075 71
rect 7165 37 7253 71
rect 7343 37 7431 71
rect 7521 37 7609 71
rect 7699 37 7787 71
rect 7877 37 7965 71
rect 8055 37 8143 71
rect 8233 37 8321 71
rect 8411 37 8499 71
rect 8589 37 8677 71
rect 8767 37 8855 71
rect -8855 -71 -8767 -37
rect -8677 -71 -8589 -37
rect -8499 -71 -8411 -37
rect -8321 -71 -8233 -37
rect -8143 -71 -8055 -37
rect -7965 -71 -7877 -37
rect -7787 -71 -7699 -37
rect -7609 -71 -7521 -37
rect -7431 -71 -7343 -37
rect -7253 -71 -7165 -37
rect -7075 -71 -6987 -37
rect -6897 -71 -6809 -37
rect -6719 -71 -6631 -37
rect -6541 -71 -6453 -37
rect -6363 -71 -6275 -37
rect -6185 -71 -6097 -37
rect -6007 -71 -5919 -37
rect -5829 -71 -5741 -37
rect -5651 -71 -5563 -37
rect -5473 -71 -5385 -37
rect -5295 -71 -5207 -37
rect -5117 -71 -5029 -37
rect -4939 -71 -4851 -37
rect -4761 -71 -4673 -37
rect -4583 -71 -4495 -37
rect -4405 -71 -4317 -37
rect -4227 -71 -4139 -37
rect -4049 -71 -3961 -37
rect -3871 -71 -3783 -37
rect -3693 -71 -3605 -37
rect -3515 -71 -3427 -37
rect -3337 -71 -3249 -37
rect -3159 -71 -3071 -37
rect -2981 -71 -2893 -37
rect -2803 -71 -2715 -37
rect -2625 -71 -2537 -37
rect -2447 -71 -2359 -37
rect -2269 -71 -2181 -37
rect -2091 -71 -2003 -37
rect -1913 -71 -1825 -37
rect -1735 -71 -1647 -37
rect -1557 -71 -1469 -37
rect -1379 -71 -1291 -37
rect -1201 -71 -1113 -37
rect -1023 -71 -935 -37
rect -845 -71 -757 -37
rect -667 -71 -579 -37
rect -489 -71 -401 -37
rect -311 -71 -223 -37
rect -133 -71 -45 -37
rect 45 -71 133 -37
rect 223 -71 311 -37
rect 401 -71 489 -37
rect 579 -71 667 -37
rect 757 -71 845 -37
rect 935 -71 1023 -37
rect 1113 -71 1201 -37
rect 1291 -71 1379 -37
rect 1469 -71 1557 -37
rect 1647 -71 1735 -37
rect 1825 -71 1913 -37
rect 2003 -71 2091 -37
rect 2181 -71 2269 -37
rect 2359 -71 2447 -37
rect 2537 -71 2625 -37
rect 2715 -71 2803 -37
rect 2893 -71 2981 -37
rect 3071 -71 3159 -37
rect 3249 -71 3337 -37
rect 3427 -71 3515 -37
rect 3605 -71 3693 -37
rect 3783 -71 3871 -37
rect 3961 -71 4049 -37
rect 4139 -71 4227 -37
rect 4317 -71 4405 -37
rect 4495 -71 4583 -37
rect 4673 -71 4761 -37
rect 4851 -71 4939 -37
rect 5029 -71 5117 -37
rect 5207 -71 5295 -37
rect 5385 -71 5473 -37
rect 5563 -71 5651 -37
rect 5741 -71 5829 -37
rect 5919 -71 6007 -37
rect 6097 -71 6185 -37
rect 6275 -71 6363 -37
rect 6453 -71 6541 -37
rect 6631 -71 6719 -37
rect 6809 -71 6897 -37
rect 6987 -71 7075 -37
rect 7165 -71 7253 -37
rect 7343 -71 7431 -37
rect 7521 -71 7609 -37
rect 7699 -71 7787 -37
rect 7877 -71 7965 -37
rect 8055 -71 8143 -37
rect 8233 -71 8321 -37
rect 8411 -71 8499 -37
rect 8589 -71 8677 -37
rect 8767 -71 8855 -37
rect -8917 -2506 -8883 -130
rect -8739 -2506 -8705 -130
rect -8561 -2506 -8527 -130
rect -8383 -2506 -8349 -130
rect -8205 -2506 -8171 -130
rect -8027 -2506 -7993 -130
rect -7849 -2506 -7815 -130
rect -7671 -2506 -7637 -130
rect -7493 -2506 -7459 -130
rect -7315 -2506 -7281 -130
rect -7137 -2506 -7103 -130
rect -6959 -2506 -6925 -130
rect -6781 -2506 -6747 -130
rect -6603 -2506 -6569 -130
rect -6425 -2506 -6391 -130
rect -6247 -2506 -6213 -130
rect -6069 -2506 -6035 -130
rect -5891 -2506 -5857 -130
rect -5713 -2506 -5679 -130
rect -5535 -2506 -5501 -130
rect -5357 -2506 -5323 -130
rect -5179 -2506 -5145 -130
rect -5001 -2506 -4967 -130
rect -4823 -2506 -4789 -130
rect -4645 -2506 -4611 -130
rect -4467 -2506 -4433 -130
rect -4289 -2506 -4255 -130
rect -4111 -2506 -4077 -130
rect -3933 -2506 -3899 -130
rect -3755 -2506 -3721 -130
rect -3577 -2506 -3543 -130
rect -3399 -2506 -3365 -130
rect -3221 -2506 -3187 -130
rect -3043 -2506 -3009 -130
rect -2865 -2506 -2831 -130
rect -2687 -2506 -2653 -130
rect -2509 -2506 -2475 -130
rect -2331 -2506 -2297 -130
rect -2153 -2506 -2119 -130
rect -1975 -2506 -1941 -130
rect -1797 -2506 -1763 -130
rect -1619 -2506 -1585 -130
rect -1441 -2506 -1407 -130
rect -1263 -2506 -1229 -130
rect -1085 -2506 -1051 -130
rect -907 -2506 -873 -130
rect -729 -2506 -695 -130
rect -551 -2506 -517 -130
rect -373 -2506 -339 -130
rect -195 -2506 -161 -130
rect -17 -2506 17 -130
rect 161 -2506 195 -130
rect 339 -2506 373 -130
rect 517 -2506 551 -130
rect 695 -2506 729 -130
rect 873 -2506 907 -130
rect 1051 -2506 1085 -130
rect 1229 -2506 1263 -130
rect 1407 -2506 1441 -130
rect 1585 -2506 1619 -130
rect 1763 -2506 1797 -130
rect 1941 -2506 1975 -130
rect 2119 -2506 2153 -130
rect 2297 -2506 2331 -130
rect 2475 -2506 2509 -130
rect 2653 -2506 2687 -130
rect 2831 -2506 2865 -130
rect 3009 -2506 3043 -130
rect 3187 -2506 3221 -130
rect 3365 -2506 3399 -130
rect 3543 -2506 3577 -130
rect 3721 -2506 3755 -130
rect 3899 -2506 3933 -130
rect 4077 -2506 4111 -130
rect 4255 -2506 4289 -130
rect 4433 -2506 4467 -130
rect 4611 -2506 4645 -130
rect 4789 -2506 4823 -130
rect 4967 -2506 5001 -130
rect 5145 -2506 5179 -130
rect 5323 -2506 5357 -130
rect 5501 -2506 5535 -130
rect 5679 -2506 5713 -130
rect 5857 -2506 5891 -130
rect 6035 -2506 6069 -130
rect 6213 -2506 6247 -130
rect 6391 -2506 6425 -130
rect 6569 -2506 6603 -130
rect 6747 -2506 6781 -130
rect 6925 -2506 6959 -130
rect 7103 -2506 7137 -130
rect 7281 -2506 7315 -130
rect 7459 -2506 7493 -130
rect 7637 -2506 7671 -130
rect 7815 -2506 7849 -130
rect 7993 -2506 8027 -130
rect 8171 -2506 8205 -130
rect 8349 -2506 8383 -130
rect 8527 -2506 8561 -130
rect 8705 -2506 8739 -130
rect 8883 -2506 8917 -130
rect -8855 -2599 -8767 -2565
rect -8677 -2599 -8589 -2565
rect -8499 -2599 -8411 -2565
rect -8321 -2599 -8233 -2565
rect -8143 -2599 -8055 -2565
rect -7965 -2599 -7877 -2565
rect -7787 -2599 -7699 -2565
rect -7609 -2599 -7521 -2565
rect -7431 -2599 -7343 -2565
rect -7253 -2599 -7165 -2565
rect -7075 -2599 -6987 -2565
rect -6897 -2599 -6809 -2565
rect -6719 -2599 -6631 -2565
rect -6541 -2599 -6453 -2565
rect -6363 -2599 -6275 -2565
rect -6185 -2599 -6097 -2565
rect -6007 -2599 -5919 -2565
rect -5829 -2599 -5741 -2565
rect -5651 -2599 -5563 -2565
rect -5473 -2599 -5385 -2565
rect -5295 -2599 -5207 -2565
rect -5117 -2599 -5029 -2565
rect -4939 -2599 -4851 -2565
rect -4761 -2599 -4673 -2565
rect -4583 -2599 -4495 -2565
rect -4405 -2599 -4317 -2565
rect -4227 -2599 -4139 -2565
rect -4049 -2599 -3961 -2565
rect -3871 -2599 -3783 -2565
rect -3693 -2599 -3605 -2565
rect -3515 -2599 -3427 -2565
rect -3337 -2599 -3249 -2565
rect -3159 -2599 -3071 -2565
rect -2981 -2599 -2893 -2565
rect -2803 -2599 -2715 -2565
rect -2625 -2599 -2537 -2565
rect -2447 -2599 -2359 -2565
rect -2269 -2599 -2181 -2565
rect -2091 -2599 -2003 -2565
rect -1913 -2599 -1825 -2565
rect -1735 -2599 -1647 -2565
rect -1557 -2599 -1469 -2565
rect -1379 -2599 -1291 -2565
rect -1201 -2599 -1113 -2565
rect -1023 -2599 -935 -2565
rect -845 -2599 -757 -2565
rect -667 -2599 -579 -2565
rect -489 -2599 -401 -2565
rect -311 -2599 -223 -2565
rect -133 -2599 -45 -2565
rect 45 -2599 133 -2565
rect 223 -2599 311 -2565
rect 401 -2599 489 -2565
rect 579 -2599 667 -2565
rect 757 -2599 845 -2565
rect 935 -2599 1023 -2565
rect 1113 -2599 1201 -2565
rect 1291 -2599 1379 -2565
rect 1469 -2599 1557 -2565
rect 1647 -2599 1735 -2565
rect 1825 -2599 1913 -2565
rect 2003 -2599 2091 -2565
rect 2181 -2599 2269 -2565
rect 2359 -2599 2447 -2565
rect 2537 -2599 2625 -2565
rect 2715 -2599 2803 -2565
rect 2893 -2599 2981 -2565
rect 3071 -2599 3159 -2565
rect 3249 -2599 3337 -2565
rect 3427 -2599 3515 -2565
rect 3605 -2599 3693 -2565
rect 3783 -2599 3871 -2565
rect 3961 -2599 4049 -2565
rect 4139 -2599 4227 -2565
rect 4317 -2599 4405 -2565
rect 4495 -2599 4583 -2565
rect 4673 -2599 4761 -2565
rect 4851 -2599 4939 -2565
rect 5029 -2599 5117 -2565
rect 5207 -2599 5295 -2565
rect 5385 -2599 5473 -2565
rect 5563 -2599 5651 -2565
rect 5741 -2599 5829 -2565
rect 5919 -2599 6007 -2565
rect 6097 -2599 6185 -2565
rect 6275 -2599 6363 -2565
rect 6453 -2599 6541 -2565
rect 6631 -2599 6719 -2565
rect 6809 -2599 6897 -2565
rect 6987 -2599 7075 -2565
rect 7165 -2599 7253 -2565
rect 7343 -2599 7431 -2565
rect 7521 -2599 7609 -2565
rect 7699 -2599 7787 -2565
rect 7877 -2599 7965 -2565
rect 8055 -2599 8143 -2565
rect 8233 -2599 8321 -2565
rect 8411 -2599 8499 -2565
rect 8589 -2599 8677 -2565
rect 8767 -2599 8855 -2565
<< metal1 >>
rect -8867 2599 -8755 2605
rect -8867 2565 -8855 2599
rect -8767 2565 -8755 2599
rect -8867 2559 -8755 2565
rect -8689 2599 -8577 2605
rect -8689 2565 -8677 2599
rect -8589 2565 -8577 2599
rect -8689 2559 -8577 2565
rect -8511 2599 -8399 2605
rect -8511 2565 -8499 2599
rect -8411 2565 -8399 2599
rect -8511 2559 -8399 2565
rect -8333 2599 -8221 2605
rect -8333 2565 -8321 2599
rect -8233 2565 -8221 2599
rect -8333 2559 -8221 2565
rect -8155 2599 -8043 2605
rect -8155 2565 -8143 2599
rect -8055 2565 -8043 2599
rect -8155 2559 -8043 2565
rect -7977 2599 -7865 2605
rect -7977 2565 -7965 2599
rect -7877 2565 -7865 2599
rect -7977 2559 -7865 2565
rect -7799 2599 -7687 2605
rect -7799 2565 -7787 2599
rect -7699 2565 -7687 2599
rect -7799 2559 -7687 2565
rect -7621 2599 -7509 2605
rect -7621 2565 -7609 2599
rect -7521 2565 -7509 2599
rect -7621 2559 -7509 2565
rect -7443 2599 -7331 2605
rect -7443 2565 -7431 2599
rect -7343 2565 -7331 2599
rect -7443 2559 -7331 2565
rect -7265 2599 -7153 2605
rect -7265 2565 -7253 2599
rect -7165 2565 -7153 2599
rect -7265 2559 -7153 2565
rect -7087 2599 -6975 2605
rect -7087 2565 -7075 2599
rect -6987 2565 -6975 2599
rect -7087 2559 -6975 2565
rect -6909 2599 -6797 2605
rect -6909 2565 -6897 2599
rect -6809 2565 -6797 2599
rect -6909 2559 -6797 2565
rect -6731 2599 -6619 2605
rect -6731 2565 -6719 2599
rect -6631 2565 -6619 2599
rect -6731 2559 -6619 2565
rect -6553 2599 -6441 2605
rect -6553 2565 -6541 2599
rect -6453 2565 -6441 2599
rect -6553 2559 -6441 2565
rect -6375 2599 -6263 2605
rect -6375 2565 -6363 2599
rect -6275 2565 -6263 2599
rect -6375 2559 -6263 2565
rect -6197 2599 -6085 2605
rect -6197 2565 -6185 2599
rect -6097 2565 -6085 2599
rect -6197 2559 -6085 2565
rect -6019 2599 -5907 2605
rect -6019 2565 -6007 2599
rect -5919 2565 -5907 2599
rect -6019 2559 -5907 2565
rect -5841 2599 -5729 2605
rect -5841 2565 -5829 2599
rect -5741 2565 -5729 2599
rect -5841 2559 -5729 2565
rect -5663 2599 -5551 2605
rect -5663 2565 -5651 2599
rect -5563 2565 -5551 2599
rect -5663 2559 -5551 2565
rect -5485 2599 -5373 2605
rect -5485 2565 -5473 2599
rect -5385 2565 -5373 2599
rect -5485 2559 -5373 2565
rect -5307 2599 -5195 2605
rect -5307 2565 -5295 2599
rect -5207 2565 -5195 2599
rect -5307 2559 -5195 2565
rect -5129 2599 -5017 2605
rect -5129 2565 -5117 2599
rect -5029 2565 -5017 2599
rect -5129 2559 -5017 2565
rect -4951 2599 -4839 2605
rect -4951 2565 -4939 2599
rect -4851 2565 -4839 2599
rect -4951 2559 -4839 2565
rect -4773 2599 -4661 2605
rect -4773 2565 -4761 2599
rect -4673 2565 -4661 2599
rect -4773 2559 -4661 2565
rect -4595 2599 -4483 2605
rect -4595 2565 -4583 2599
rect -4495 2565 -4483 2599
rect -4595 2559 -4483 2565
rect -4417 2599 -4305 2605
rect -4417 2565 -4405 2599
rect -4317 2565 -4305 2599
rect -4417 2559 -4305 2565
rect -4239 2599 -4127 2605
rect -4239 2565 -4227 2599
rect -4139 2565 -4127 2599
rect -4239 2559 -4127 2565
rect -4061 2599 -3949 2605
rect -4061 2565 -4049 2599
rect -3961 2565 -3949 2599
rect -4061 2559 -3949 2565
rect -3883 2599 -3771 2605
rect -3883 2565 -3871 2599
rect -3783 2565 -3771 2599
rect -3883 2559 -3771 2565
rect -3705 2599 -3593 2605
rect -3705 2565 -3693 2599
rect -3605 2565 -3593 2599
rect -3705 2559 -3593 2565
rect -3527 2599 -3415 2605
rect -3527 2565 -3515 2599
rect -3427 2565 -3415 2599
rect -3527 2559 -3415 2565
rect -3349 2599 -3237 2605
rect -3349 2565 -3337 2599
rect -3249 2565 -3237 2599
rect -3349 2559 -3237 2565
rect -3171 2599 -3059 2605
rect -3171 2565 -3159 2599
rect -3071 2565 -3059 2599
rect -3171 2559 -3059 2565
rect -2993 2599 -2881 2605
rect -2993 2565 -2981 2599
rect -2893 2565 -2881 2599
rect -2993 2559 -2881 2565
rect -2815 2599 -2703 2605
rect -2815 2565 -2803 2599
rect -2715 2565 -2703 2599
rect -2815 2559 -2703 2565
rect -2637 2599 -2525 2605
rect -2637 2565 -2625 2599
rect -2537 2565 -2525 2599
rect -2637 2559 -2525 2565
rect -2459 2599 -2347 2605
rect -2459 2565 -2447 2599
rect -2359 2565 -2347 2599
rect -2459 2559 -2347 2565
rect -2281 2599 -2169 2605
rect -2281 2565 -2269 2599
rect -2181 2565 -2169 2599
rect -2281 2559 -2169 2565
rect -2103 2599 -1991 2605
rect -2103 2565 -2091 2599
rect -2003 2565 -1991 2599
rect -2103 2559 -1991 2565
rect -1925 2599 -1813 2605
rect -1925 2565 -1913 2599
rect -1825 2565 -1813 2599
rect -1925 2559 -1813 2565
rect -1747 2599 -1635 2605
rect -1747 2565 -1735 2599
rect -1647 2565 -1635 2599
rect -1747 2559 -1635 2565
rect -1569 2599 -1457 2605
rect -1569 2565 -1557 2599
rect -1469 2565 -1457 2599
rect -1569 2559 -1457 2565
rect -1391 2599 -1279 2605
rect -1391 2565 -1379 2599
rect -1291 2565 -1279 2599
rect -1391 2559 -1279 2565
rect -1213 2599 -1101 2605
rect -1213 2565 -1201 2599
rect -1113 2565 -1101 2599
rect -1213 2559 -1101 2565
rect -1035 2599 -923 2605
rect -1035 2565 -1023 2599
rect -935 2565 -923 2599
rect -1035 2559 -923 2565
rect -857 2599 -745 2605
rect -857 2565 -845 2599
rect -757 2565 -745 2599
rect -857 2559 -745 2565
rect -679 2599 -567 2605
rect -679 2565 -667 2599
rect -579 2565 -567 2599
rect -679 2559 -567 2565
rect -501 2599 -389 2605
rect -501 2565 -489 2599
rect -401 2565 -389 2599
rect -501 2559 -389 2565
rect -323 2599 -211 2605
rect -323 2565 -311 2599
rect -223 2565 -211 2599
rect -323 2559 -211 2565
rect -145 2599 -33 2605
rect -145 2565 -133 2599
rect -45 2565 -33 2599
rect -145 2559 -33 2565
rect 33 2599 145 2605
rect 33 2565 45 2599
rect 133 2565 145 2599
rect 33 2559 145 2565
rect 211 2599 323 2605
rect 211 2565 223 2599
rect 311 2565 323 2599
rect 211 2559 323 2565
rect 389 2599 501 2605
rect 389 2565 401 2599
rect 489 2565 501 2599
rect 389 2559 501 2565
rect 567 2599 679 2605
rect 567 2565 579 2599
rect 667 2565 679 2599
rect 567 2559 679 2565
rect 745 2599 857 2605
rect 745 2565 757 2599
rect 845 2565 857 2599
rect 745 2559 857 2565
rect 923 2599 1035 2605
rect 923 2565 935 2599
rect 1023 2565 1035 2599
rect 923 2559 1035 2565
rect 1101 2599 1213 2605
rect 1101 2565 1113 2599
rect 1201 2565 1213 2599
rect 1101 2559 1213 2565
rect 1279 2599 1391 2605
rect 1279 2565 1291 2599
rect 1379 2565 1391 2599
rect 1279 2559 1391 2565
rect 1457 2599 1569 2605
rect 1457 2565 1469 2599
rect 1557 2565 1569 2599
rect 1457 2559 1569 2565
rect 1635 2599 1747 2605
rect 1635 2565 1647 2599
rect 1735 2565 1747 2599
rect 1635 2559 1747 2565
rect 1813 2599 1925 2605
rect 1813 2565 1825 2599
rect 1913 2565 1925 2599
rect 1813 2559 1925 2565
rect 1991 2599 2103 2605
rect 1991 2565 2003 2599
rect 2091 2565 2103 2599
rect 1991 2559 2103 2565
rect 2169 2599 2281 2605
rect 2169 2565 2181 2599
rect 2269 2565 2281 2599
rect 2169 2559 2281 2565
rect 2347 2599 2459 2605
rect 2347 2565 2359 2599
rect 2447 2565 2459 2599
rect 2347 2559 2459 2565
rect 2525 2599 2637 2605
rect 2525 2565 2537 2599
rect 2625 2565 2637 2599
rect 2525 2559 2637 2565
rect 2703 2599 2815 2605
rect 2703 2565 2715 2599
rect 2803 2565 2815 2599
rect 2703 2559 2815 2565
rect 2881 2599 2993 2605
rect 2881 2565 2893 2599
rect 2981 2565 2993 2599
rect 2881 2559 2993 2565
rect 3059 2599 3171 2605
rect 3059 2565 3071 2599
rect 3159 2565 3171 2599
rect 3059 2559 3171 2565
rect 3237 2599 3349 2605
rect 3237 2565 3249 2599
rect 3337 2565 3349 2599
rect 3237 2559 3349 2565
rect 3415 2599 3527 2605
rect 3415 2565 3427 2599
rect 3515 2565 3527 2599
rect 3415 2559 3527 2565
rect 3593 2599 3705 2605
rect 3593 2565 3605 2599
rect 3693 2565 3705 2599
rect 3593 2559 3705 2565
rect 3771 2599 3883 2605
rect 3771 2565 3783 2599
rect 3871 2565 3883 2599
rect 3771 2559 3883 2565
rect 3949 2599 4061 2605
rect 3949 2565 3961 2599
rect 4049 2565 4061 2599
rect 3949 2559 4061 2565
rect 4127 2599 4239 2605
rect 4127 2565 4139 2599
rect 4227 2565 4239 2599
rect 4127 2559 4239 2565
rect 4305 2599 4417 2605
rect 4305 2565 4317 2599
rect 4405 2565 4417 2599
rect 4305 2559 4417 2565
rect 4483 2599 4595 2605
rect 4483 2565 4495 2599
rect 4583 2565 4595 2599
rect 4483 2559 4595 2565
rect 4661 2599 4773 2605
rect 4661 2565 4673 2599
rect 4761 2565 4773 2599
rect 4661 2559 4773 2565
rect 4839 2599 4951 2605
rect 4839 2565 4851 2599
rect 4939 2565 4951 2599
rect 4839 2559 4951 2565
rect 5017 2599 5129 2605
rect 5017 2565 5029 2599
rect 5117 2565 5129 2599
rect 5017 2559 5129 2565
rect 5195 2599 5307 2605
rect 5195 2565 5207 2599
rect 5295 2565 5307 2599
rect 5195 2559 5307 2565
rect 5373 2599 5485 2605
rect 5373 2565 5385 2599
rect 5473 2565 5485 2599
rect 5373 2559 5485 2565
rect 5551 2599 5663 2605
rect 5551 2565 5563 2599
rect 5651 2565 5663 2599
rect 5551 2559 5663 2565
rect 5729 2599 5841 2605
rect 5729 2565 5741 2599
rect 5829 2565 5841 2599
rect 5729 2559 5841 2565
rect 5907 2599 6019 2605
rect 5907 2565 5919 2599
rect 6007 2565 6019 2599
rect 5907 2559 6019 2565
rect 6085 2599 6197 2605
rect 6085 2565 6097 2599
rect 6185 2565 6197 2599
rect 6085 2559 6197 2565
rect 6263 2599 6375 2605
rect 6263 2565 6275 2599
rect 6363 2565 6375 2599
rect 6263 2559 6375 2565
rect 6441 2599 6553 2605
rect 6441 2565 6453 2599
rect 6541 2565 6553 2599
rect 6441 2559 6553 2565
rect 6619 2599 6731 2605
rect 6619 2565 6631 2599
rect 6719 2565 6731 2599
rect 6619 2559 6731 2565
rect 6797 2599 6909 2605
rect 6797 2565 6809 2599
rect 6897 2565 6909 2599
rect 6797 2559 6909 2565
rect 6975 2599 7087 2605
rect 6975 2565 6987 2599
rect 7075 2565 7087 2599
rect 6975 2559 7087 2565
rect 7153 2599 7265 2605
rect 7153 2565 7165 2599
rect 7253 2565 7265 2599
rect 7153 2559 7265 2565
rect 7331 2599 7443 2605
rect 7331 2565 7343 2599
rect 7431 2565 7443 2599
rect 7331 2559 7443 2565
rect 7509 2599 7621 2605
rect 7509 2565 7521 2599
rect 7609 2565 7621 2599
rect 7509 2559 7621 2565
rect 7687 2599 7799 2605
rect 7687 2565 7699 2599
rect 7787 2565 7799 2599
rect 7687 2559 7799 2565
rect 7865 2599 7977 2605
rect 7865 2565 7877 2599
rect 7965 2565 7977 2599
rect 7865 2559 7977 2565
rect 8043 2599 8155 2605
rect 8043 2565 8055 2599
rect 8143 2565 8155 2599
rect 8043 2559 8155 2565
rect 8221 2599 8333 2605
rect 8221 2565 8233 2599
rect 8321 2565 8333 2599
rect 8221 2559 8333 2565
rect 8399 2599 8511 2605
rect 8399 2565 8411 2599
rect 8499 2565 8511 2599
rect 8399 2559 8511 2565
rect 8577 2599 8689 2605
rect 8577 2565 8589 2599
rect 8677 2565 8689 2599
rect 8577 2559 8689 2565
rect 8755 2599 8867 2605
rect 8755 2565 8767 2599
rect 8855 2565 8867 2599
rect 8755 2559 8867 2565
rect -8923 2506 -8877 2518
rect -8923 130 -8917 2506
rect -8883 130 -8877 2506
rect -8923 118 -8877 130
rect -8745 2506 -8699 2518
rect -8745 130 -8739 2506
rect -8705 130 -8699 2506
rect -8745 118 -8699 130
rect -8567 2506 -8521 2518
rect -8567 130 -8561 2506
rect -8527 130 -8521 2506
rect -8567 118 -8521 130
rect -8389 2506 -8343 2518
rect -8389 130 -8383 2506
rect -8349 130 -8343 2506
rect -8389 118 -8343 130
rect -8211 2506 -8165 2518
rect -8211 130 -8205 2506
rect -8171 130 -8165 2506
rect -8211 118 -8165 130
rect -8033 2506 -7987 2518
rect -8033 130 -8027 2506
rect -7993 130 -7987 2506
rect -8033 118 -7987 130
rect -7855 2506 -7809 2518
rect -7855 130 -7849 2506
rect -7815 130 -7809 2506
rect -7855 118 -7809 130
rect -7677 2506 -7631 2518
rect -7677 130 -7671 2506
rect -7637 130 -7631 2506
rect -7677 118 -7631 130
rect -7499 2506 -7453 2518
rect -7499 130 -7493 2506
rect -7459 130 -7453 2506
rect -7499 118 -7453 130
rect -7321 2506 -7275 2518
rect -7321 130 -7315 2506
rect -7281 130 -7275 2506
rect -7321 118 -7275 130
rect -7143 2506 -7097 2518
rect -7143 130 -7137 2506
rect -7103 130 -7097 2506
rect -7143 118 -7097 130
rect -6965 2506 -6919 2518
rect -6965 130 -6959 2506
rect -6925 130 -6919 2506
rect -6965 118 -6919 130
rect -6787 2506 -6741 2518
rect -6787 130 -6781 2506
rect -6747 130 -6741 2506
rect -6787 118 -6741 130
rect -6609 2506 -6563 2518
rect -6609 130 -6603 2506
rect -6569 130 -6563 2506
rect -6609 118 -6563 130
rect -6431 2506 -6385 2518
rect -6431 130 -6425 2506
rect -6391 130 -6385 2506
rect -6431 118 -6385 130
rect -6253 2506 -6207 2518
rect -6253 130 -6247 2506
rect -6213 130 -6207 2506
rect -6253 118 -6207 130
rect -6075 2506 -6029 2518
rect -6075 130 -6069 2506
rect -6035 130 -6029 2506
rect -6075 118 -6029 130
rect -5897 2506 -5851 2518
rect -5897 130 -5891 2506
rect -5857 130 -5851 2506
rect -5897 118 -5851 130
rect -5719 2506 -5673 2518
rect -5719 130 -5713 2506
rect -5679 130 -5673 2506
rect -5719 118 -5673 130
rect -5541 2506 -5495 2518
rect -5541 130 -5535 2506
rect -5501 130 -5495 2506
rect -5541 118 -5495 130
rect -5363 2506 -5317 2518
rect -5363 130 -5357 2506
rect -5323 130 -5317 2506
rect -5363 118 -5317 130
rect -5185 2506 -5139 2518
rect -5185 130 -5179 2506
rect -5145 130 -5139 2506
rect -5185 118 -5139 130
rect -5007 2506 -4961 2518
rect -5007 130 -5001 2506
rect -4967 130 -4961 2506
rect -5007 118 -4961 130
rect -4829 2506 -4783 2518
rect -4829 130 -4823 2506
rect -4789 130 -4783 2506
rect -4829 118 -4783 130
rect -4651 2506 -4605 2518
rect -4651 130 -4645 2506
rect -4611 130 -4605 2506
rect -4651 118 -4605 130
rect -4473 2506 -4427 2518
rect -4473 130 -4467 2506
rect -4433 130 -4427 2506
rect -4473 118 -4427 130
rect -4295 2506 -4249 2518
rect -4295 130 -4289 2506
rect -4255 130 -4249 2506
rect -4295 118 -4249 130
rect -4117 2506 -4071 2518
rect -4117 130 -4111 2506
rect -4077 130 -4071 2506
rect -4117 118 -4071 130
rect -3939 2506 -3893 2518
rect -3939 130 -3933 2506
rect -3899 130 -3893 2506
rect -3939 118 -3893 130
rect -3761 2506 -3715 2518
rect -3761 130 -3755 2506
rect -3721 130 -3715 2506
rect -3761 118 -3715 130
rect -3583 2506 -3537 2518
rect -3583 130 -3577 2506
rect -3543 130 -3537 2506
rect -3583 118 -3537 130
rect -3405 2506 -3359 2518
rect -3405 130 -3399 2506
rect -3365 130 -3359 2506
rect -3405 118 -3359 130
rect -3227 2506 -3181 2518
rect -3227 130 -3221 2506
rect -3187 130 -3181 2506
rect -3227 118 -3181 130
rect -3049 2506 -3003 2518
rect -3049 130 -3043 2506
rect -3009 130 -3003 2506
rect -3049 118 -3003 130
rect -2871 2506 -2825 2518
rect -2871 130 -2865 2506
rect -2831 130 -2825 2506
rect -2871 118 -2825 130
rect -2693 2506 -2647 2518
rect -2693 130 -2687 2506
rect -2653 130 -2647 2506
rect -2693 118 -2647 130
rect -2515 2506 -2469 2518
rect -2515 130 -2509 2506
rect -2475 130 -2469 2506
rect -2515 118 -2469 130
rect -2337 2506 -2291 2518
rect -2337 130 -2331 2506
rect -2297 130 -2291 2506
rect -2337 118 -2291 130
rect -2159 2506 -2113 2518
rect -2159 130 -2153 2506
rect -2119 130 -2113 2506
rect -2159 118 -2113 130
rect -1981 2506 -1935 2518
rect -1981 130 -1975 2506
rect -1941 130 -1935 2506
rect -1981 118 -1935 130
rect -1803 2506 -1757 2518
rect -1803 130 -1797 2506
rect -1763 130 -1757 2506
rect -1803 118 -1757 130
rect -1625 2506 -1579 2518
rect -1625 130 -1619 2506
rect -1585 130 -1579 2506
rect -1625 118 -1579 130
rect -1447 2506 -1401 2518
rect -1447 130 -1441 2506
rect -1407 130 -1401 2506
rect -1447 118 -1401 130
rect -1269 2506 -1223 2518
rect -1269 130 -1263 2506
rect -1229 130 -1223 2506
rect -1269 118 -1223 130
rect -1091 2506 -1045 2518
rect -1091 130 -1085 2506
rect -1051 130 -1045 2506
rect -1091 118 -1045 130
rect -913 2506 -867 2518
rect -913 130 -907 2506
rect -873 130 -867 2506
rect -913 118 -867 130
rect -735 2506 -689 2518
rect -735 130 -729 2506
rect -695 130 -689 2506
rect -735 118 -689 130
rect -557 2506 -511 2518
rect -557 130 -551 2506
rect -517 130 -511 2506
rect -557 118 -511 130
rect -379 2506 -333 2518
rect -379 130 -373 2506
rect -339 130 -333 2506
rect -379 118 -333 130
rect -201 2506 -155 2518
rect -201 130 -195 2506
rect -161 130 -155 2506
rect -201 118 -155 130
rect -23 2506 23 2518
rect -23 130 -17 2506
rect 17 130 23 2506
rect -23 118 23 130
rect 155 2506 201 2518
rect 155 130 161 2506
rect 195 130 201 2506
rect 155 118 201 130
rect 333 2506 379 2518
rect 333 130 339 2506
rect 373 130 379 2506
rect 333 118 379 130
rect 511 2506 557 2518
rect 511 130 517 2506
rect 551 130 557 2506
rect 511 118 557 130
rect 689 2506 735 2518
rect 689 130 695 2506
rect 729 130 735 2506
rect 689 118 735 130
rect 867 2506 913 2518
rect 867 130 873 2506
rect 907 130 913 2506
rect 867 118 913 130
rect 1045 2506 1091 2518
rect 1045 130 1051 2506
rect 1085 130 1091 2506
rect 1045 118 1091 130
rect 1223 2506 1269 2518
rect 1223 130 1229 2506
rect 1263 130 1269 2506
rect 1223 118 1269 130
rect 1401 2506 1447 2518
rect 1401 130 1407 2506
rect 1441 130 1447 2506
rect 1401 118 1447 130
rect 1579 2506 1625 2518
rect 1579 130 1585 2506
rect 1619 130 1625 2506
rect 1579 118 1625 130
rect 1757 2506 1803 2518
rect 1757 130 1763 2506
rect 1797 130 1803 2506
rect 1757 118 1803 130
rect 1935 2506 1981 2518
rect 1935 130 1941 2506
rect 1975 130 1981 2506
rect 1935 118 1981 130
rect 2113 2506 2159 2518
rect 2113 130 2119 2506
rect 2153 130 2159 2506
rect 2113 118 2159 130
rect 2291 2506 2337 2518
rect 2291 130 2297 2506
rect 2331 130 2337 2506
rect 2291 118 2337 130
rect 2469 2506 2515 2518
rect 2469 130 2475 2506
rect 2509 130 2515 2506
rect 2469 118 2515 130
rect 2647 2506 2693 2518
rect 2647 130 2653 2506
rect 2687 130 2693 2506
rect 2647 118 2693 130
rect 2825 2506 2871 2518
rect 2825 130 2831 2506
rect 2865 130 2871 2506
rect 2825 118 2871 130
rect 3003 2506 3049 2518
rect 3003 130 3009 2506
rect 3043 130 3049 2506
rect 3003 118 3049 130
rect 3181 2506 3227 2518
rect 3181 130 3187 2506
rect 3221 130 3227 2506
rect 3181 118 3227 130
rect 3359 2506 3405 2518
rect 3359 130 3365 2506
rect 3399 130 3405 2506
rect 3359 118 3405 130
rect 3537 2506 3583 2518
rect 3537 130 3543 2506
rect 3577 130 3583 2506
rect 3537 118 3583 130
rect 3715 2506 3761 2518
rect 3715 130 3721 2506
rect 3755 130 3761 2506
rect 3715 118 3761 130
rect 3893 2506 3939 2518
rect 3893 130 3899 2506
rect 3933 130 3939 2506
rect 3893 118 3939 130
rect 4071 2506 4117 2518
rect 4071 130 4077 2506
rect 4111 130 4117 2506
rect 4071 118 4117 130
rect 4249 2506 4295 2518
rect 4249 130 4255 2506
rect 4289 130 4295 2506
rect 4249 118 4295 130
rect 4427 2506 4473 2518
rect 4427 130 4433 2506
rect 4467 130 4473 2506
rect 4427 118 4473 130
rect 4605 2506 4651 2518
rect 4605 130 4611 2506
rect 4645 130 4651 2506
rect 4605 118 4651 130
rect 4783 2506 4829 2518
rect 4783 130 4789 2506
rect 4823 130 4829 2506
rect 4783 118 4829 130
rect 4961 2506 5007 2518
rect 4961 130 4967 2506
rect 5001 130 5007 2506
rect 4961 118 5007 130
rect 5139 2506 5185 2518
rect 5139 130 5145 2506
rect 5179 130 5185 2506
rect 5139 118 5185 130
rect 5317 2506 5363 2518
rect 5317 130 5323 2506
rect 5357 130 5363 2506
rect 5317 118 5363 130
rect 5495 2506 5541 2518
rect 5495 130 5501 2506
rect 5535 130 5541 2506
rect 5495 118 5541 130
rect 5673 2506 5719 2518
rect 5673 130 5679 2506
rect 5713 130 5719 2506
rect 5673 118 5719 130
rect 5851 2506 5897 2518
rect 5851 130 5857 2506
rect 5891 130 5897 2506
rect 5851 118 5897 130
rect 6029 2506 6075 2518
rect 6029 130 6035 2506
rect 6069 130 6075 2506
rect 6029 118 6075 130
rect 6207 2506 6253 2518
rect 6207 130 6213 2506
rect 6247 130 6253 2506
rect 6207 118 6253 130
rect 6385 2506 6431 2518
rect 6385 130 6391 2506
rect 6425 130 6431 2506
rect 6385 118 6431 130
rect 6563 2506 6609 2518
rect 6563 130 6569 2506
rect 6603 130 6609 2506
rect 6563 118 6609 130
rect 6741 2506 6787 2518
rect 6741 130 6747 2506
rect 6781 130 6787 2506
rect 6741 118 6787 130
rect 6919 2506 6965 2518
rect 6919 130 6925 2506
rect 6959 130 6965 2506
rect 6919 118 6965 130
rect 7097 2506 7143 2518
rect 7097 130 7103 2506
rect 7137 130 7143 2506
rect 7097 118 7143 130
rect 7275 2506 7321 2518
rect 7275 130 7281 2506
rect 7315 130 7321 2506
rect 7275 118 7321 130
rect 7453 2506 7499 2518
rect 7453 130 7459 2506
rect 7493 130 7499 2506
rect 7453 118 7499 130
rect 7631 2506 7677 2518
rect 7631 130 7637 2506
rect 7671 130 7677 2506
rect 7631 118 7677 130
rect 7809 2506 7855 2518
rect 7809 130 7815 2506
rect 7849 130 7855 2506
rect 7809 118 7855 130
rect 7987 2506 8033 2518
rect 7987 130 7993 2506
rect 8027 130 8033 2506
rect 7987 118 8033 130
rect 8165 2506 8211 2518
rect 8165 130 8171 2506
rect 8205 130 8211 2506
rect 8165 118 8211 130
rect 8343 2506 8389 2518
rect 8343 130 8349 2506
rect 8383 130 8389 2506
rect 8343 118 8389 130
rect 8521 2506 8567 2518
rect 8521 130 8527 2506
rect 8561 130 8567 2506
rect 8521 118 8567 130
rect 8699 2506 8745 2518
rect 8699 130 8705 2506
rect 8739 130 8745 2506
rect 8699 118 8745 130
rect 8877 2506 8923 2518
rect 8877 130 8883 2506
rect 8917 130 8923 2506
rect 8877 118 8923 130
rect -8867 71 -8755 77
rect -8867 37 -8855 71
rect -8767 37 -8755 71
rect -8867 31 -8755 37
rect -8689 71 -8577 77
rect -8689 37 -8677 71
rect -8589 37 -8577 71
rect -8689 31 -8577 37
rect -8511 71 -8399 77
rect -8511 37 -8499 71
rect -8411 37 -8399 71
rect -8511 31 -8399 37
rect -8333 71 -8221 77
rect -8333 37 -8321 71
rect -8233 37 -8221 71
rect -8333 31 -8221 37
rect -8155 71 -8043 77
rect -8155 37 -8143 71
rect -8055 37 -8043 71
rect -8155 31 -8043 37
rect -7977 71 -7865 77
rect -7977 37 -7965 71
rect -7877 37 -7865 71
rect -7977 31 -7865 37
rect -7799 71 -7687 77
rect -7799 37 -7787 71
rect -7699 37 -7687 71
rect -7799 31 -7687 37
rect -7621 71 -7509 77
rect -7621 37 -7609 71
rect -7521 37 -7509 71
rect -7621 31 -7509 37
rect -7443 71 -7331 77
rect -7443 37 -7431 71
rect -7343 37 -7331 71
rect -7443 31 -7331 37
rect -7265 71 -7153 77
rect -7265 37 -7253 71
rect -7165 37 -7153 71
rect -7265 31 -7153 37
rect -7087 71 -6975 77
rect -7087 37 -7075 71
rect -6987 37 -6975 71
rect -7087 31 -6975 37
rect -6909 71 -6797 77
rect -6909 37 -6897 71
rect -6809 37 -6797 71
rect -6909 31 -6797 37
rect -6731 71 -6619 77
rect -6731 37 -6719 71
rect -6631 37 -6619 71
rect -6731 31 -6619 37
rect -6553 71 -6441 77
rect -6553 37 -6541 71
rect -6453 37 -6441 71
rect -6553 31 -6441 37
rect -6375 71 -6263 77
rect -6375 37 -6363 71
rect -6275 37 -6263 71
rect -6375 31 -6263 37
rect -6197 71 -6085 77
rect -6197 37 -6185 71
rect -6097 37 -6085 71
rect -6197 31 -6085 37
rect -6019 71 -5907 77
rect -6019 37 -6007 71
rect -5919 37 -5907 71
rect -6019 31 -5907 37
rect -5841 71 -5729 77
rect -5841 37 -5829 71
rect -5741 37 -5729 71
rect -5841 31 -5729 37
rect -5663 71 -5551 77
rect -5663 37 -5651 71
rect -5563 37 -5551 71
rect -5663 31 -5551 37
rect -5485 71 -5373 77
rect -5485 37 -5473 71
rect -5385 37 -5373 71
rect -5485 31 -5373 37
rect -5307 71 -5195 77
rect -5307 37 -5295 71
rect -5207 37 -5195 71
rect -5307 31 -5195 37
rect -5129 71 -5017 77
rect -5129 37 -5117 71
rect -5029 37 -5017 71
rect -5129 31 -5017 37
rect -4951 71 -4839 77
rect -4951 37 -4939 71
rect -4851 37 -4839 71
rect -4951 31 -4839 37
rect -4773 71 -4661 77
rect -4773 37 -4761 71
rect -4673 37 -4661 71
rect -4773 31 -4661 37
rect -4595 71 -4483 77
rect -4595 37 -4583 71
rect -4495 37 -4483 71
rect -4595 31 -4483 37
rect -4417 71 -4305 77
rect -4417 37 -4405 71
rect -4317 37 -4305 71
rect -4417 31 -4305 37
rect -4239 71 -4127 77
rect -4239 37 -4227 71
rect -4139 37 -4127 71
rect -4239 31 -4127 37
rect -4061 71 -3949 77
rect -4061 37 -4049 71
rect -3961 37 -3949 71
rect -4061 31 -3949 37
rect -3883 71 -3771 77
rect -3883 37 -3871 71
rect -3783 37 -3771 71
rect -3883 31 -3771 37
rect -3705 71 -3593 77
rect -3705 37 -3693 71
rect -3605 37 -3593 71
rect -3705 31 -3593 37
rect -3527 71 -3415 77
rect -3527 37 -3515 71
rect -3427 37 -3415 71
rect -3527 31 -3415 37
rect -3349 71 -3237 77
rect -3349 37 -3337 71
rect -3249 37 -3237 71
rect -3349 31 -3237 37
rect -3171 71 -3059 77
rect -3171 37 -3159 71
rect -3071 37 -3059 71
rect -3171 31 -3059 37
rect -2993 71 -2881 77
rect -2993 37 -2981 71
rect -2893 37 -2881 71
rect -2993 31 -2881 37
rect -2815 71 -2703 77
rect -2815 37 -2803 71
rect -2715 37 -2703 71
rect -2815 31 -2703 37
rect -2637 71 -2525 77
rect -2637 37 -2625 71
rect -2537 37 -2525 71
rect -2637 31 -2525 37
rect -2459 71 -2347 77
rect -2459 37 -2447 71
rect -2359 37 -2347 71
rect -2459 31 -2347 37
rect -2281 71 -2169 77
rect -2281 37 -2269 71
rect -2181 37 -2169 71
rect -2281 31 -2169 37
rect -2103 71 -1991 77
rect -2103 37 -2091 71
rect -2003 37 -1991 71
rect -2103 31 -1991 37
rect -1925 71 -1813 77
rect -1925 37 -1913 71
rect -1825 37 -1813 71
rect -1925 31 -1813 37
rect -1747 71 -1635 77
rect -1747 37 -1735 71
rect -1647 37 -1635 71
rect -1747 31 -1635 37
rect -1569 71 -1457 77
rect -1569 37 -1557 71
rect -1469 37 -1457 71
rect -1569 31 -1457 37
rect -1391 71 -1279 77
rect -1391 37 -1379 71
rect -1291 37 -1279 71
rect -1391 31 -1279 37
rect -1213 71 -1101 77
rect -1213 37 -1201 71
rect -1113 37 -1101 71
rect -1213 31 -1101 37
rect -1035 71 -923 77
rect -1035 37 -1023 71
rect -935 37 -923 71
rect -1035 31 -923 37
rect -857 71 -745 77
rect -857 37 -845 71
rect -757 37 -745 71
rect -857 31 -745 37
rect -679 71 -567 77
rect -679 37 -667 71
rect -579 37 -567 71
rect -679 31 -567 37
rect -501 71 -389 77
rect -501 37 -489 71
rect -401 37 -389 71
rect -501 31 -389 37
rect -323 71 -211 77
rect -323 37 -311 71
rect -223 37 -211 71
rect -323 31 -211 37
rect -145 71 -33 77
rect -145 37 -133 71
rect -45 37 -33 71
rect -145 31 -33 37
rect 33 71 145 77
rect 33 37 45 71
rect 133 37 145 71
rect 33 31 145 37
rect 211 71 323 77
rect 211 37 223 71
rect 311 37 323 71
rect 211 31 323 37
rect 389 71 501 77
rect 389 37 401 71
rect 489 37 501 71
rect 389 31 501 37
rect 567 71 679 77
rect 567 37 579 71
rect 667 37 679 71
rect 567 31 679 37
rect 745 71 857 77
rect 745 37 757 71
rect 845 37 857 71
rect 745 31 857 37
rect 923 71 1035 77
rect 923 37 935 71
rect 1023 37 1035 71
rect 923 31 1035 37
rect 1101 71 1213 77
rect 1101 37 1113 71
rect 1201 37 1213 71
rect 1101 31 1213 37
rect 1279 71 1391 77
rect 1279 37 1291 71
rect 1379 37 1391 71
rect 1279 31 1391 37
rect 1457 71 1569 77
rect 1457 37 1469 71
rect 1557 37 1569 71
rect 1457 31 1569 37
rect 1635 71 1747 77
rect 1635 37 1647 71
rect 1735 37 1747 71
rect 1635 31 1747 37
rect 1813 71 1925 77
rect 1813 37 1825 71
rect 1913 37 1925 71
rect 1813 31 1925 37
rect 1991 71 2103 77
rect 1991 37 2003 71
rect 2091 37 2103 71
rect 1991 31 2103 37
rect 2169 71 2281 77
rect 2169 37 2181 71
rect 2269 37 2281 71
rect 2169 31 2281 37
rect 2347 71 2459 77
rect 2347 37 2359 71
rect 2447 37 2459 71
rect 2347 31 2459 37
rect 2525 71 2637 77
rect 2525 37 2537 71
rect 2625 37 2637 71
rect 2525 31 2637 37
rect 2703 71 2815 77
rect 2703 37 2715 71
rect 2803 37 2815 71
rect 2703 31 2815 37
rect 2881 71 2993 77
rect 2881 37 2893 71
rect 2981 37 2993 71
rect 2881 31 2993 37
rect 3059 71 3171 77
rect 3059 37 3071 71
rect 3159 37 3171 71
rect 3059 31 3171 37
rect 3237 71 3349 77
rect 3237 37 3249 71
rect 3337 37 3349 71
rect 3237 31 3349 37
rect 3415 71 3527 77
rect 3415 37 3427 71
rect 3515 37 3527 71
rect 3415 31 3527 37
rect 3593 71 3705 77
rect 3593 37 3605 71
rect 3693 37 3705 71
rect 3593 31 3705 37
rect 3771 71 3883 77
rect 3771 37 3783 71
rect 3871 37 3883 71
rect 3771 31 3883 37
rect 3949 71 4061 77
rect 3949 37 3961 71
rect 4049 37 4061 71
rect 3949 31 4061 37
rect 4127 71 4239 77
rect 4127 37 4139 71
rect 4227 37 4239 71
rect 4127 31 4239 37
rect 4305 71 4417 77
rect 4305 37 4317 71
rect 4405 37 4417 71
rect 4305 31 4417 37
rect 4483 71 4595 77
rect 4483 37 4495 71
rect 4583 37 4595 71
rect 4483 31 4595 37
rect 4661 71 4773 77
rect 4661 37 4673 71
rect 4761 37 4773 71
rect 4661 31 4773 37
rect 4839 71 4951 77
rect 4839 37 4851 71
rect 4939 37 4951 71
rect 4839 31 4951 37
rect 5017 71 5129 77
rect 5017 37 5029 71
rect 5117 37 5129 71
rect 5017 31 5129 37
rect 5195 71 5307 77
rect 5195 37 5207 71
rect 5295 37 5307 71
rect 5195 31 5307 37
rect 5373 71 5485 77
rect 5373 37 5385 71
rect 5473 37 5485 71
rect 5373 31 5485 37
rect 5551 71 5663 77
rect 5551 37 5563 71
rect 5651 37 5663 71
rect 5551 31 5663 37
rect 5729 71 5841 77
rect 5729 37 5741 71
rect 5829 37 5841 71
rect 5729 31 5841 37
rect 5907 71 6019 77
rect 5907 37 5919 71
rect 6007 37 6019 71
rect 5907 31 6019 37
rect 6085 71 6197 77
rect 6085 37 6097 71
rect 6185 37 6197 71
rect 6085 31 6197 37
rect 6263 71 6375 77
rect 6263 37 6275 71
rect 6363 37 6375 71
rect 6263 31 6375 37
rect 6441 71 6553 77
rect 6441 37 6453 71
rect 6541 37 6553 71
rect 6441 31 6553 37
rect 6619 71 6731 77
rect 6619 37 6631 71
rect 6719 37 6731 71
rect 6619 31 6731 37
rect 6797 71 6909 77
rect 6797 37 6809 71
rect 6897 37 6909 71
rect 6797 31 6909 37
rect 6975 71 7087 77
rect 6975 37 6987 71
rect 7075 37 7087 71
rect 6975 31 7087 37
rect 7153 71 7265 77
rect 7153 37 7165 71
rect 7253 37 7265 71
rect 7153 31 7265 37
rect 7331 71 7443 77
rect 7331 37 7343 71
rect 7431 37 7443 71
rect 7331 31 7443 37
rect 7509 71 7621 77
rect 7509 37 7521 71
rect 7609 37 7621 71
rect 7509 31 7621 37
rect 7687 71 7799 77
rect 7687 37 7699 71
rect 7787 37 7799 71
rect 7687 31 7799 37
rect 7865 71 7977 77
rect 7865 37 7877 71
rect 7965 37 7977 71
rect 7865 31 7977 37
rect 8043 71 8155 77
rect 8043 37 8055 71
rect 8143 37 8155 71
rect 8043 31 8155 37
rect 8221 71 8333 77
rect 8221 37 8233 71
rect 8321 37 8333 71
rect 8221 31 8333 37
rect 8399 71 8511 77
rect 8399 37 8411 71
rect 8499 37 8511 71
rect 8399 31 8511 37
rect 8577 71 8689 77
rect 8577 37 8589 71
rect 8677 37 8689 71
rect 8577 31 8689 37
rect 8755 71 8867 77
rect 8755 37 8767 71
rect 8855 37 8867 71
rect 8755 31 8867 37
rect -8867 -37 -8755 -31
rect -8867 -71 -8855 -37
rect -8767 -71 -8755 -37
rect -8867 -77 -8755 -71
rect -8689 -37 -8577 -31
rect -8689 -71 -8677 -37
rect -8589 -71 -8577 -37
rect -8689 -77 -8577 -71
rect -8511 -37 -8399 -31
rect -8511 -71 -8499 -37
rect -8411 -71 -8399 -37
rect -8511 -77 -8399 -71
rect -8333 -37 -8221 -31
rect -8333 -71 -8321 -37
rect -8233 -71 -8221 -37
rect -8333 -77 -8221 -71
rect -8155 -37 -8043 -31
rect -8155 -71 -8143 -37
rect -8055 -71 -8043 -37
rect -8155 -77 -8043 -71
rect -7977 -37 -7865 -31
rect -7977 -71 -7965 -37
rect -7877 -71 -7865 -37
rect -7977 -77 -7865 -71
rect -7799 -37 -7687 -31
rect -7799 -71 -7787 -37
rect -7699 -71 -7687 -37
rect -7799 -77 -7687 -71
rect -7621 -37 -7509 -31
rect -7621 -71 -7609 -37
rect -7521 -71 -7509 -37
rect -7621 -77 -7509 -71
rect -7443 -37 -7331 -31
rect -7443 -71 -7431 -37
rect -7343 -71 -7331 -37
rect -7443 -77 -7331 -71
rect -7265 -37 -7153 -31
rect -7265 -71 -7253 -37
rect -7165 -71 -7153 -37
rect -7265 -77 -7153 -71
rect -7087 -37 -6975 -31
rect -7087 -71 -7075 -37
rect -6987 -71 -6975 -37
rect -7087 -77 -6975 -71
rect -6909 -37 -6797 -31
rect -6909 -71 -6897 -37
rect -6809 -71 -6797 -37
rect -6909 -77 -6797 -71
rect -6731 -37 -6619 -31
rect -6731 -71 -6719 -37
rect -6631 -71 -6619 -37
rect -6731 -77 -6619 -71
rect -6553 -37 -6441 -31
rect -6553 -71 -6541 -37
rect -6453 -71 -6441 -37
rect -6553 -77 -6441 -71
rect -6375 -37 -6263 -31
rect -6375 -71 -6363 -37
rect -6275 -71 -6263 -37
rect -6375 -77 -6263 -71
rect -6197 -37 -6085 -31
rect -6197 -71 -6185 -37
rect -6097 -71 -6085 -37
rect -6197 -77 -6085 -71
rect -6019 -37 -5907 -31
rect -6019 -71 -6007 -37
rect -5919 -71 -5907 -37
rect -6019 -77 -5907 -71
rect -5841 -37 -5729 -31
rect -5841 -71 -5829 -37
rect -5741 -71 -5729 -37
rect -5841 -77 -5729 -71
rect -5663 -37 -5551 -31
rect -5663 -71 -5651 -37
rect -5563 -71 -5551 -37
rect -5663 -77 -5551 -71
rect -5485 -37 -5373 -31
rect -5485 -71 -5473 -37
rect -5385 -71 -5373 -37
rect -5485 -77 -5373 -71
rect -5307 -37 -5195 -31
rect -5307 -71 -5295 -37
rect -5207 -71 -5195 -37
rect -5307 -77 -5195 -71
rect -5129 -37 -5017 -31
rect -5129 -71 -5117 -37
rect -5029 -71 -5017 -37
rect -5129 -77 -5017 -71
rect -4951 -37 -4839 -31
rect -4951 -71 -4939 -37
rect -4851 -71 -4839 -37
rect -4951 -77 -4839 -71
rect -4773 -37 -4661 -31
rect -4773 -71 -4761 -37
rect -4673 -71 -4661 -37
rect -4773 -77 -4661 -71
rect -4595 -37 -4483 -31
rect -4595 -71 -4583 -37
rect -4495 -71 -4483 -37
rect -4595 -77 -4483 -71
rect -4417 -37 -4305 -31
rect -4417 -71 -4405 -37
rect -4317 -71 -4305 -37
rect -4417 -77 -4305 -71
rect -4239 -37 -4127 -31
rect -4239 -71 -4227 -37
rect -4139 -71 -4127 -37
rect -4239 -77 -4127 -71
rect -4061 -37 -3949 -31
rect -4061 -71 -4049 -37
rect -3961 -71 -3949 -37
rect -4061 -77 -3949 -71
rect -3883 -37 -3771 -31
rect -3883 -71 -3871 -37
rect -3783 -71 -3771 -37
rect -3883 -77 -3771 -71
rect -3705 -37 -3593 -31
rect -3705 -71 -3693 -37
rect -3605 -71 -3593 -37
rect -3705 -77 -3593 -71
rect -3527 -37 -3415 -31
rect -3527 -71 -3515 -37
rect -3427 -71 -3415 -37
rect -3527 -77 -3415 -71
rect -3349 -37 -3237 -31
rect -3349 -71 -3337 -37
rect -3249 -71 -3237 -37
rect -3349 -77 -3237 -71
rect -3171 -37 -3059 -31
rect -3171 -71 -3159 -37
rect -3071 -71 -3059 -37
rect -3171 -77 -3059 -71
rect -2993 -37 -2881 -31
rect -2993 -71 -2981 -37
rect -2893 -71 -2881 -37
rect -2993 -77 -2881 -71
rect -2815 -37 -2703 -31
rect -2815 -71 -2803 -37
rect -2715 -71 -2703 -37
rect -2815 -77 -2703 -71
rect -2637 -37 -2525 -31
rect -2637 -71 -2625 -37
rect -2537 -71 -2525 -37
rect -2637 -77 -2525 -71
rect -2459 -37 -2347 -31
rect -2459 -71 -2447 -37
rect -2359 -71 -2347 -37
rect -2459 -77 -2347 -71
rect -2281 -37 -2169 -31
rect -2281 -71 -2269 -37
rect -2181 -71 -2169 -37
rect -2281 -77 -2169 -71
rect -2103 -37 -1991 -31
rect -2103 -71 -2091 -37
rect -2003 -71 -1991 -37
rect -2103 -77 -1991 -71
rect -1925 -37 -1813 -31
rect -1925 -71 -1913 -37
rect -1825 -71 -1813 -37
rect -1925 -77 -1813 -71
rect -1747 -37 -1635 -31
rect -1747 -71 -1735 -37
rect -1647 -71 -1635 -37
rect -1747 -77 -1635 -71
rect -1569 -37 -1457 -31
rect -1569 -71 -1557 -37
rect -1469 -71 -1457 -37
rect -1569 -77 -1457 -71
rect -1391 -37 -1279 -31
rect -1391 -71 -1379 -37
rect -1291 -71 -1279 -37
rect -1391 -77 -1279 -71
rect -1213 -37 -1101 -31
rect -1213 -71 -1201 -37
rect -1113 -71 -1101 -37
rect -1213 -77 -1101 -71
rect -1035 -37 -923 -31
rect -1035 -71 -1023 -37
rect -935 -71 -923 -37
rect -1035 -77 -923 -71
rect -857 -37 -745 -31
rect -857 -71 -845 -37
rect -757 -71 -745 -37
rect -857 -77 -745 -71
rect -679 -37 -567 -31
rect -679 -71 -667 -37
rect -579 -71 -567 -37
rect -679 -77 -567 -71
rect -501 -37 -389 -31
rect -501 -71 -489 -37
rect -401 -71 -389 -37
rect -501 -77 -389 -71
rect -323 -37 -211 -31
rect -323 -71 -311 -37
rect -223 -71 -211 -37
rect -323 -77 -211 -71
rect -145 -37 -33 -31
rect -145 -71 -133 -37
rect -45 -71 -33 -37
rect -145 -77 -33 -71
rect 33 -37 145 -31
rect 33 -71 45 -37
rect 133 -71 145 -37
rect 33 -77 145 -71
rect 211 -37 323 -31
rect 211 -71 223 -37
rect 311 -71 323 -37
rect 211 -77 323 -71
rect 389 -37 501 -31
rect 389 -71 401 -37
rect 489 -71 501 -37
rect 389 -77 501 -71
rect 567 -37 679 -31
rect 567 -71 579 -37
rect 667 -71 679 -37
rect 567 -77 679 -71
rect 745 -37 857 -31
rect 745 -71 757 -37
rect 845 -71 857 -37
rect 745 -77 857 -71
rect 923 -37 1035 -31
rect 923 -71 935 -37
rect 1023 -71 1035 -37
rect 923 -77 1035 -71
rect 1101 -37 1213 -31
rect 1101 -71 1113 -37
rect 1201 -71 1213 -37
rect 1101 -77 1213 -71
rect 1279 -37 1391 -31
rect 1279 -71 1291 -37
rect 1379 -71 1391 -37
rect 1279 -77 1391 -71
rect 1457 -37 1569 -31
rect 1457 -71 1469 -37
rect 1557 -71 1569 -37
rect 1457 -77 1569 -71
rect 1635 -37 1747 -31
rect 1635 -71 1647 -37
rect 1735 -71 1747 -37
rect 1635 -77 1747 -71
rect 1813 -37 1925 -31
rect 1813 -71 1825 -37
rect 1913 -71 1925 -37
rect 1813 -77 1925 -71
rect 1991 -37 2103 -31
rect 1991 -71 2003 -37
rect 2091 -71 2103 -37
rect 1991 -77 2103 -71
rect 2169 -37 2281 -31
rect 2169 -71 2181 -37
rect 2269 -71 2281 -37
rect 2169 -77 2281 -71
rect 2347 -37 2459 -31
rect 2347 -71 2359 -37
rect 2447 -71 2459 -37
rect 2347 -77 2459 -71
rect 2525 -37 2637 -31
rect 2525 -71 2537 -37
rect 2625 -71 2637 -37
rect 2525 -77 2637 -71
rect 2703 -37 2815 -31
rect 2703 -71 2715 -37
rect 2803 -71 2815 -37
rect 2703 -77 2815 -71
rect 2881 -37 2993 -31
rect 2881 -71 2893 -37
rect 2981 -71 2993 -37
rect 2881 -77 2993 -71
rect 3059 -37 3171 -31
rect 3059 -71 3071 -37
rect 3159 -71 3171 -37
rect 3059 -77 3171 -71
rect 3237 -37 3349 -31
rect 3237 -71 3249 -37
rect 3337 -71 3349 -37
rect 3237 -77 3349 -71
rect 3415 -37 3527 -31
rect 3415 -71 3427 -37
rect 3515 -71 3527 -37
rect 3415 -77 3527 -71
rect 3593 -37 3705 -31
rect 3593 -71 3605 -37
rect 3693 -71 3705 -37
rect 3593 -77 3705 -71
rect 3771 -37 3883 -31
rect 3771 -71 3783 -37
rect 3871 -71 3883 -37
rect 3771 -77 3883 -71
rect 3949 -37 4061 -31
rect 3949 -71 3961 -37
rect 4049 -71 4061 -37
rect 3949 -77 4061 -71
rect 4127 -37 4239 -31
rect 4127 -71 4139 -37
rect 4227 -71 4239 -37
rect 4127 -77 4239 -71
rect 4305 -37 4417 -31
rect 4305 -71 4317 -37
rect 4405 -71 4417 -37
rect 4305 -77 4417 -71
rect 4483 -37 4595 -31
rect 4483 -71 4495 -37
rect 4583 -71 4595 -37
rect 4483 -77 4595 -71
rect 4661 -37 4773 -31
rect 4661 -71 4673 -37
rect 4761 -71 4773 -37
rect 4661 -77 4773 -71
rect 4839 -37 4951 -31
rect 4839 -71 4851 -37
rect 4939 -71 4951 -37
rect 4839 -77 4951 -71
rect 5017 -37 5129 -31
rect 5017 -71 5029 -37
rect 5117 -71 5129 -37
rect 5017 -77 5129 -71
rect 5195 -37 5307 -31
rect 5195 -71 5207 -37
rect 5295 -71 5307 -37
rect 5195 -77 5307 -71
rect 5373 -37 5485 -31
rect 5373 -71 5385 -37
rect 5473 -71 5485 -37
rect 5373 -77 5485 -71
rect 5551 -37 5663 -31
rect 5551 -71 5563 -37
rect 5651 -71 5663 -37
rect 5551 -77 5663 -71
rect 5729 -37 5841 -31
rect 5729 -71 5741 -37
rect 5829 -71 5841 -37
rect 5729 -77 5841 -71
rect 5907 -37 6019 -31
rect 5907 -71 5919 -37
rect 6007 -71 6019 -37
rect 5907 -77 6019 -71
rect 6085 -37 6197 -31
rect 6085 -71 6097 -37
rect 6185 -71 6197 -37
rect 6085 -77 6197 -71
rect 6263 -37 6375 -31
rect 6263 -71 6275 -37
rect 6363 -71 6375 -37
rect 6263 -77 6375 -71
rect 6441 -37 6553 -31
rect 6441 -71 6453 -37
rect 6541 -71 6553 -37
rect 6441 -77 6553 -71
rect 6619 -37 6731 -31
rect 6619 -71 6631 -37
rect 6719 -71 6731 -37
rect 6619 -77 6731 -71
rect 6797 -37 6909 -31
rect 6797 -71 6809 -37
rect 6897 -71 6909 -37
rect 6797 -77 6909 -71
rect 6975 -37 7087 -31
rect 6975 -71 6987 -37
rect 7075 -71 7087 -37
rect 6975 -77 7087 -71
rect 7153 -37 7265 -31
rect 7153 -71 7165 -37
rect 7253 -71 7265 -37
rect 7153 -77 7265 -71
rect 7331 -37 7443 -31
rect 7331 -71 7343 -37
rect 7431 -71 7443 -37
rect 7331 -77 7443 -71
rect 7509 -37 7621 -31
rect 7509 -71 7521 -37
rect 7609 -71 7621 -37
rect 7509 -77 7621 -71
rect 7687 -37 7799 -31
rect 7687 -71 7699 -37
rect 7787 -71 7799 -37
rect 7687 -77 7799 -71
rect 7865 -37 7977 -31
rect 7865 -71 7877 -37
rect 7965 -71 7977 -37
rect 7865 -77 7977 -71
rect 8043 -37 8155 -31
rect 8043 -71 8055 -37
rect 8143 -71 8155 -37
rect 8043 -77 8155 -71
rect 8221 -37 8333 -31
rect 8221 -71 8233 -37
rect 8321 -71 8333 -37
rect 8221 -77 8333 -71
rect 8399 -37 8511 -31
rect 8399 -71 8411 -37
rect 8499 -71 8511 -37
rect 8399 -77 8511 -71
rect 8577 -37 8689 -31
rect 8577 -71 8589 -37
rect 8677 -71 8689 -37
rect 8577 -77 8689 -71
rect 8755 -37 8867 -31
rect 8755 -71 8767 -37
rect 8855 -71 8867 -37
rect 8755 -77 8867 -71
rect -8923 -130 -8877 -118
rect -8923 -2506 -8917 -130
rect -8883 -2506 -8877 -130
rect -8923 -2518 -8877 -2506
rect -8745 -130 -8699 -118
rect -8745 -2506 -8739 -130
rect -8705 -2506 -8699 -130
rect -8745 -2518 -8699 -2506
rect -8567 -130 -8521 -118
rect -8567 -2506 -8561 -130
rect -8527 -2506 -8521 -130
rect -8567 -2518 -8521 -2506
rect -8389 -130 -8343 -118
rect -8389 -2506 -8383 -130
rect -8349 -2506 -8343 -130
rect -8389 -2518 -8343 -2506
rect -8211 -130 -8165 -118
rect -8211 -2506 -8205 -130
rect -8171 -2506 -8165 -130
rect -8211 -2518 -8165 -2506
rect -8033 -130 -7987 -118
rect -8033 -2506 -8027 -130
rect -7993 -2506 -7987 -130
rect -8033 -2518 -7987 -2506
rect -7855 -130 -7809 -118
rect -7855 -2506 -7849 -130
rect -7815 -2506 -7809 -130
rect -7855 -2518 -7809 -2506
rect -7677 -130 -7631 -118
rect -7677 -2506 -7671 -130
rect -7637 -2506 -7631 -130
rect -7677 -2518 -7631 -2506
rect -7499 -130 -7453 -118
rect -7499 -2506 -7493 -130
rect -7459 -2506 -7453 -130
rect -7499 -2518 -7453 -2506
rect -7321 -130 -7275 -118
rect -7321 -2506 -7315 -130
rect -7281 -2506 -7275 -130
rect -7321 -2518 -7275 -2506
rect -7143 -130 -7097 -118
rect -7143 -2506 -7137 -130
rect -7103 -2506 -7097 -130
rect -7143 -2518 -7097 -2506
rect -6965 -130 -6919 -118
rect -6965 -2506 -6959 -130
rect -6925 -2506 -6919 -130
rect -6965 -2518 -6919 -2506
rect -6787 -130 -6741 -118
rect -6787 -2506 -6781 -130
rect -6747 -2506 -6741 -130
rect -6787 -2518 -6741 -2506
rect -6609 -130 -6563 -118
rect -6609 -2506 -6603 -130
rect -6569 -2506 -6563 -130
rect -6609 -2518 -6563 -2506
rect -6431 -130 -6385 -118
rect -6431 -2506 -6425 -130
rect -6391 -2506 -6385 -130
rect -6431 -2518 -6385 -2506
rect -6253 -130 -6207 -118
rect -6253 -2506 -6247 -130
rect -6213 -2506 -6207 -130
rect -6253 -2518 -6207 -2506
rect -6075 -130 -6029 -118
rect -6075 -2506 -6069 -130
rect -6035 -2506 -6029 -130
rect -6075 -2518 -6029 -2506
rect -5897 -130 -5851 -118
rect -5897 -2506 -5891 -130
rect -5857 -2506 -5851 -130
rect -5897 -2518 -5851 -2506
rect -5719 -130 -5673 -118
rect -5719 -2506 -5713 -130
rect -5679 -2506 -5673 -130
rect -5719 -2518 -5673 -2506
rect -5541 -130 -5495 -118
rect -5541 -2506 -5535 -130
rect -5501 -2506 -5495 -130
rect -5541 -2518 -5495 -2506
rect -5363 -130 -5317 -118
rect -5363 -2506 -5357 -130
rect -5323 -2506 -5317 -130
rect -5363 -2518 -5317 -2506
rect -5185 -130 -5139 -118
rect -5185 -2506 -5179 -130
rect -5145 -2506 -5139 -130
rect -5185 -2518 -5139 -2506
rect -5007 -130 -4961 -118
rect -5007 -2506 -5001 -130
rect -4967 -2506 -4961 -130
rect -5007 -2518 -4961 -2506
rect -4829 -130 -4783 -118
rect -4829 -2506 -4823 -130
rect -4789 -2506 -4783 -130
rect -4829 -2518 -4783 -2506
rect -4651 -130 -4605 -118
rect -4651 -2506 -4645 -130
rect -4611 -2506 -4605 -130
rect -4651 -2518 -4605 -2506
rect -4473 -130 -4427 -118
rect -4473 -2506 -4467 -130
rect -4433 -2506 -4427 -130
rect -4473 -2518 -4427 -2506
rect -4295 -130 -4249 -118
rect -4295 -2506 -4289 -130
rect -4255 -2506 -4249 -130
rect -4295 -2518 -4249 -2506
rect -4117 -130 -4071 -118
rect -4117 -2506 -4111 -130
rect -4077 -2506 -4071 -130
rect -4117 -2518 -4071 -2506
rect -3939 -130 -3893 -118
rect -3939 -2506 -3933 -130
rect -3899 -2506 -3893 -130
rect -3939 -2518 -3893 -2506
rect -3761 -130 -3715 -118
rect -3761 -2506 -3755 -130
rect -3721 -2506 -3715 -130
rect -3761 -2518 -3715 -2506
rect -3583 -130 -3537 -118
rect -3583 -2506 -3577 -130
rect -3543 -2506 -3537 -130
rect -3583 -2518 -3537 -2506
rect -3405 -130 -3359 -118
rect -3405 -2506 -3399 -130
rect -3365 -2506 -3359 -130
rect -3405 -2518 -3359 -2506
rect -3227 -130 -3181 -118
rect -3227 -2506 -3221 -130
rect -3187 -2506 -3181 -130
rect -3227 -2518 -3181 -2506
rect -3049 -130 -3003 -118
rect -3049 -2506 -3043 -130
rect -3009 -2506 -3003 -130
rect -3049 -2518 -3003 -2506
rect -2871 -130 -2825 -118
rect -2871 -2506 -2865 -130
rect -2831 -2506 -2825 -130
rect -2871 -2518 -2825 -2506
rect -2693 -130 -2647 -118
rect -2693 -2506 -2687 -130
rect -2653 -2506 -2647 -130
rect -2693 -2518 -2647 -2506
rect -2515 -130 -2469 -118
rect -2515 -2506 -2509 -130
rect -2475 -2506 -2469 -130
rect -2515 -2518 -2469 -2506
rect -2337 -130 -2291 -118
rect -2337 -2506 -2331 -130
rect -2297 -2506 -2291 -130
rect -2337 -2518 -2291 -2506
rect -2159 -130 -2113 -118
rect -2159 -2506 -2153 -130
rect -2119 -2506 -2113 -130
rect -2159 -2518 -2113 -2506
rect -1981 -130 -1935 -118
rect -1981 -2506 -1975 -130
rect -1941 -2506 -1935 -130
rect -1981 -2518 -1935 -2506
rect -1803 -130 -1757 -118
rect -1803 -2506 -1797 -130
rect -1763 -2506 -1757 -130
rect -1803 -2518 -1757 -2506
rect -1625 -130 -1579 -118
rect -1625 -2506 -1619 -130
rect -1585 -2506 -1579 -130
rect -1625 -2518 -1579 -2506
rect -1447 -130 -1401 -118
rect -1447 -2506 -1441 -130
rect -1407 -2506 -1401 -130
rect -1447 -2518 -1401 -2506
rect -1269 -130 -1223 -118
rect -1269 -2506 -1263 -130
rect -1229 -2506 -1223 -130
rect -1269 -2518 -1223 -2506
rect -1091 -130 -1045 -118
rect -1091 -2506 -1085 -130
rect -1051 -2506 -1045 -130
rect -1091 -2518 -1045 -2506
rect -913 -130 -867 -118
rect -913 -2506 -907 -130
rect -873 -2506 -867 -130
rect -913 -2518 -867 -2506
rect -735 -130 -689 -118
rect -735 -2506 -729 -130
rect -695 -2506 -689 -130
rect -735 -2518 -689 -2506
rect -557 -130 -511 -118
rect -557 -2506 -551 -130
rect -517 -2506 -511 -130
rect -557 -2518 -511 -2506
rect -379 -130 -333 -118
rect -379 -2506 -373 -130
rect -339 -2506 -333 -130
rect -379 -2518 -333 -2506
rect -201 -130 -155 -118
rect -201 -2506 -195 -130
rect -161 -2506 -155 -130
rect -201 -2518 -155 -2506
rect -23 -130 23 -118
rect -23 -2506 -17 -130
rect 17 -2506 23 -130
rect -23 -2518 23 -2506
rect 155 -130 201 -118
rect 155 -2506 161 -130
rect 195 -2506 201 -130
rect 155 -2518 201 -2506
rect 333 -130 379 -118
rect 333 -2506 339 -130
rect 373 -2506 379 -130
rect 333 -2518 379 -2506
rect 511 -130 557 -118
rect 511 -2506 517 -130
rect 551 -2506 557 -130
rect 511 -2518 557 -2506
rect 689 -130 735 -118
rect 689 -2506 695 -130
rect 729 -2506 735 -130
rect 689 -2518 735 -2506
rect 867 -130 913 -118
rect 867 -2506 873 -130
rect 907 -2506 913 -130
rect 867 -2518 913 -2506
rect 1045 -130 1091 -118
rect 1045 -2506 1051 -130
rect 1085 -2506 1091 -130
rect 1045 -2518 1091 -2506
rect 1223 -130 1269 -118
rect 1223 -2506 1229 -130
rect 1263 -2506 1269 -130
rect 1223 -2518 1269 -2506
rect 1401 -130 1447 -118
rect 1401 -2506 1407 -130
rect 1441 -2506 1447 -130
rect 1401 -2518 1447 -2506
rect 1579 -130 1625 -118
rect 1579 -2506 1585 -130
rect 1619 -2506 1625 -130
rect 1579 -2518 1625 -2506
rect 1757 -130 1803 -118
rect 1757 -2506 1763 -130
rect 1797 -2506 1803 -130
rect 1757 -2518 1803 -2506
rect 1935 -130 1981 -118
rect 1935 -2506 1941 -130
rect 1975 -2506 1981 -130
rect 1935 -2518 1981 -2506
rect 2113 -130 2159 -118
rect 2113 -2506 2119 -130
rect 2153 -2506 2159 -130
rect 2113 -2518 2159 -2506
rect 2291 -130 2337 -118
rect 2291 -2506 2297 -130
rect 2331 -2506 2337 -130
rect 2291 -2518 2337 -2506
rect 2469 -130 2515 -118
rect 2469 -2506 2475 -130
rect 2509 -2506 2515 -130
rect 2469 -2518 2515 -2506
rect 2647 -130 2693 -118
rect 2647 -2506 2653 -130
rect 2687 -2506 2693 -130
rect 2647 -2518 2693 -2506
rect 2825 -130 2871 -118
rect 2825 -2506 2831 -130
rect 2865 -2506 2871 -130
rect 2825 -2518 2871 -2506
rect 3003 -130 3049 -118
rect 3003 -2506 3009 -130
rect 3043 -2506 3049 -130
rect 3003 -2518 3049 -2506
rect 3181 -130 3227 -118
rect 3181 -2506 3187 -130
rect 3221 -2506 3227 -130
rect 3181 -2518 3227 -2506
rect 3359 -130 3405 -118
rect 3359 -2506 3365 -130
rect 3399 -2506 3405 -130
rect 3359 -2518 3405 -2506
rect 3537 -130 3583 -118
rect 3537 -2506 3543 -130
rect 3577 -2506 3583 -130
rect 3537 -2518 3583 -2506
rect 3715 -130 3761 -118
rect 3715 -2506 3721 -130
rect 3755 -2506 3761 -130
rect 3715 -2518 3761 -2506
rect 3893 -130 3939 -118
rect 3893 -2506 3899 -130
rect 3933 -2506 3939 -130
rect 3893 -2518 3939 -2506
rect 4071 -130 4117 -118
rect 4071 -2506 4077 -130
rect 4111 -2506 4117 -130
rect 4071 -2518 4117 -2506
rect 4249 -130 4295 -118
rect 4249 -2506 4255 -130
rect 4289 -2506 4295 -130
rect 4249 -2518 4295 -2506
rect 4427 -130 4473 -118
rect 4427 -2506 4433 -130
rect 4467 -2506 4473 -130
rect 4427 -2518 4473 -2506
rect 4605 -130 4651 -118
rect 4605 -2506 4611 -130
rect 4645 -2506 4651 -130
rect 4605 -2518 4651 -2506
rect 4783 -130 4829 -118
rect 4783 -2506 4789 -130
rect 4823 -2506 4829 -130
rect 4783 -2518 4829 -2506
rect 4961 -130 5007 -118
rect 4961 -2506 4967 -130
rect 5001 -2506 5007 -130
rect 4961 -2518 5007 -2506
rect 5139 -130 5185 -118
rect 5139 -2506 5145 -130
rect 5179 -2506 5185 -130
rect 5139 -2518 5185 -2506
rect 5317 -130 5363 -118
rect 5317 -2506 5323 -130
rect 5357 -2506 5363 -130
rect 5317 -2518 5363 -2506
rect 5495 -130 5541 -118
rect 5495 -2506 5501 -130
rect 5535 -2506 5541 -130
rect 5495 -2518 5541 -2506
rect 5673 -130 5719 -118
rect 5673 -2506 5679 -130
rect 5713 -2506 5719 -130
rect 5673 -2518 5719 -2506
rect 5851 -130 5897 -118
rect 5851 -2506 5857 -130
rect 5891 -2506 5897 -130
rect 5851 -2518 5897 -2506
rect 6029 -130 6075 -118
rect 6029 -2506 6035 -130
rect 6069 -2506 6075 -130
rect 6029 -2518 6075 -2506
rect 6207 -130 6253 -118
rect 6207 -2506 6213 -130
rect 6247 -2506 6253 -130
rect 6207 -2518 6253 -2506
rect 6385 -130 6431 -118
rect 6385 -2506 6391 -130
rect 6425 -2506 6431 -130
rect 6385 -2518 6431 -2506
rect 6563 -130 6609 -118
rect 6563 -2506 6569 -130
rect 6603 -2506 6609 -130
rect 6563 -2518 6609 -2506
rect 6741 -130 6787 -118
rect 6741 -2506 6747 -130
rect 6781 -2506 6787 -130
rect 6741 -2518 6787 -2506
rect 6919 -130 6965 -118
rect 6919 -2506 6925 -130
rect 6959 -2506 6965 -130
rect 6919 -2518 6965 -2506
rect 7097 -130 7143 -118
rect 7097 -2506 7103 -130
rect 7137 -2506 7143 -130
rect 7097 -2518 7143 -2506
rect 7275 -130 7321 -118
rect 7275 -2506 7281 -130
rect 7315 -2506 7321 -130
rect 7275 -2518 7321 -2506
rect 7453 -130 7499 -118
rect 7453 -2506 7459 -130
rect 7493 -2506 7499 -130
rect 7453 -2518 7499 -2506
rect 7631 -130 7677 -118
rect 7631 -2506 7637 -130
rect 7671 -2506 7677 -130
rect 7631 -2518 7677 -2506
rect 7809 -130 7855 -118
rect 7809 -2506 7815 -130
rect 7849 -2506 7855 -130
rect 7809 -2518 7855 -2506
rect 7987 -130 8033 -118
rect 7987 -2506 7993 -130
rect 8027 -2506 8033 -130
rect 7987 -2518 8033 -2506
rect 8165 -130 8211 -118
rect 8165 -2506 8171 -130
rect 8205 -2506 8211 -130
rect 8165 -2518 8211 -2506
rect 8343 -130 8389 -118
rect 8343 -2506 8349 -130
rect 8383 -2506 8389 -130
rect 8343 -2518 8389 -2506
rect 8521 -130 8567 -118
rect 8521 -2506 8527 -130
rect 8561 -2506 8567 -130
rect 8521 -2518 8567 -2506
rect 8699 -130 8745 -118
rect 8699 -2506 8705 -130
rect 8739 -2506 8745 -130
rect 8699 -2518 8745 -2506
rect 8877 -130 8923 -118
rect 8877 -2506 8883 -130
rect 8917 -2506 8923 -130
rect 8877 -2518 8923 -2506
rect -8867 -2565 -8755 -2559
rect -8867 -2599 -8855 -2565
rect -8767 -2599 -8755 -2565
rect -8867 -2605 -8755 -2599
rect -8689 -2565 -8577 -2559
rect -8689 -2599 -8677 -2565
rect -8589 -2599 -8577 -2565
rect -8689 -2605 -8577 -2599
rect -8511 -2565 -8399 -2559
rect -8511 -2599 -8499 -2565
rect -8411 -2599 -8399 -2565
rect -8511 -2605 -8399 -2599
rect -8333 -2565 -8221 -2559
rect -8333 -2599 -8321 -2565
rect -8233 -2599 -8221 -2565
rect -8333 -2605 -8221 -2599
rect -8155 -2565 -8043 -2559
rect -8155 -2599 -8143 -2565
rect -8055 -2599 -8043 -2565
rect -8155 -2605 -8043 -2599
rect -7977 -2565 -7865 -2559
rect -7977 -2599 -7965 -2565
rect -7877 -2599 -7865 -2565
rect -7977 -2605 -7865 -2599
rect -7799 -2565 -7687 -2559
rect -7799 -2599 -7787 -2565
rect -7699 -2599 -7687 -2565
rect -7799 -2605 -7687 -2599
rect -7621 -2565 -7509 -2559
rect -7621 -2599 -7609 -2565
rect -7521 -2599 -7509 -2565
rect -7621 -2605 -7509 -2599
rect -7443 -2565 -7331 -2559
rect -7443 -2599 -7431 -2565
rect -7343 -2599 -7331 -2565
rect -7443 -2605 -7331 -2599
rect -7265 -2565 -7153 -2559
rect -7265 -2599 -7253 -2565
rect -7165 -2599 -7153 -2565
rect -7265 -2605 -7153 -2599
rect -7087 -2565 -6975 -2559
rect -7087 -2599 -7075 -2565
rect -6987 -2599 -6975 -2565
rect -7087 -2605 -6975 -2599
rect -6909 -2565 -6797 -2559
rect -6909 -2599 -6897 -2565
rect -6809 -2599 -6797 -2565
rect -6909 -2605 -6797 -2599
rect -6731 -2565 -6619 -2559
rect -6731 -2599 -6719 -2565
rect -6631 -2599 -6619 -2565
rect -6731 -2605 -6619 -2599
rect -6553 -2565 -6441 -2559
rect -6553 -2599 -6541 -2565
rect -6453 -2599 -6441 -2565
rect -6553 -2605 -6441 -2599
rect -6375 -2565 -6263 -2559
rect -6375 -2599 -6363 -2565
rect -6275 -2599 -6263 -2565
rect -6375 -2605 -6263 -2599
rect -6197 -2565 -6085 -2559
rect -6197 -2599 -6185 -2565
rect -6097 -2599 -6085 -2565
rect -6197 -2605 -6085 -2599
rect -6019 -2565 -5907 -2559
rect -6019 -2599 -6007 -2565
rect -5919 -2599 -5907 -2565
rect -6019 -2605 -5907 -2599
rect -5841 -2565 -5729 -2559
rect -5841 -2599 -5829 -2565
rect -5741 -2599 -5729 -2565
rect -5841 -2605 -5729 -2599
rect -5663 -2565 -5551 -2559
rect -5663 -2599 -5651 -2565
rect -5563 -2599 -5551 -2565
rect -5663 -2605 -5551 -2599
rect -5485 -2565 -5373 -2559
rect -5485 -2599 -5473 -2565
rect -5385 -2599 -5373 -2565
rect -5485 -2605 -5373 -2599
rect -5307 -2565 -5195 -2559
rect -5307 -2599 -5295 -2565
rect -5207 -2599 -5195 -2565
rect -5307 -2605 -5195 -2599
rect -5129 -2565 -5017 -2559
rect -5129 -2599 -5117 -2565
rect -5029 -2599 -5017 -2565
rect -5129 -2605 -5017 -2599
rect -4951 -2565 -4839 -2559
rect -4951 -2599 -4939 -2565
rect -4851 -2599 -4839 -2565
rect -4951 -2605 -4839 -2599
rect -4773 -2565 -4661 -2559
rect -4773 -2599 -4761 -2565
rect -4673 -2599 -4661 -2565
rect -4773 -2605 -4661 -2599
rect -4595 -2565 -4483 -2559
rect -4595 -2599 -4583 -2565
rect -4495 -2599 -4483 -2565
rect -4595 -2605 -4483 -2599
rect -4417 -2565 -4305 -2559
rect -4417 -2599 -4405 -2565
rect -4317 -2599 -4305 -2565
rect -4417 -2605 -4305 -2599
rect -4239 -2565 -4127 -2559
rect -4239 -2599 -4227 -2565
rect -4139 -2599 -4127 -2565
rect -4239 -2605 -4127 -2599
rect -4061 -2565 -3949 -2559
rect -4061 -2599 -4049 -2565
rect -3961 -2599 -3949 -2565
rect -4061 -2605 -3949 -2599
rect -3883 -2565 -3771 -2559
rect -3883 -2599 -3871 -2565
rect -3783 -2599 -3771 -2565
rect -3883 -2605 -3771 -2599
rect -3705 -2565 -3593 -2559
rect -3705 -2599 -3693 -2565
rect -3605 -2599 -3593 -2565
rect -3705 -2605 -3593 -2599
rect -3527 -2565 -3415 -2559
rect -3527 -2599 -3515 -2565
rect -3427 -2599 -3415 -2565
rect -3527 -2605 -3415 -2599
rect -3349 -2565 -3237 -2559
rect -3349 -2599 -3337 -2565
rect -3249 -2599 -3237 -2565
rect -3349 -2605 -3237 -2599
rect -3171 -2565 -3059 -2559
rect -3171 -2599 -3159 -2565
rect -3071 -2599 -3059 -2565
rect -3171 -2605 -3059 -2599
rect -2993 -2565 -2881 -2559
rect -2993 -2599 -2981 -2565
rect -2893 -2599 -2881 -2565
rect -2993 -2605 -2881 -2599
rect -2815 -2565 -2703 -2559
rect -2815 -2599 -2803 -2565
rect -2715 -2599 -2703 -2565
rect -2815 -2605 -2703 -2599
rect -2637 -2565 -2525 -2559
rect -2637 -2599 -2625 -2565
rect -2537 -2599 -2525 -2565
rect -2637 -2605 -2525 -2599
rect -2459 -2565 -2347 -2559
rect -2459 -2599 -2447 -2565
rect -2359 -2599 -2347 -2565
rect -2459 -2605 -2347 -2599
rect -2281 -2565 -2169 -2559
rect -2281 -2599 -2269 -2565
rect -2181 -2599 -2169 -2565
rect -2281 -2605 -2169 -2599
rect -2103 -2565 -1991 -2559
rect -2103 -2599 -2091 -2565
rect -2003 -2599 -1991 -2565
rect -2103 -2605 -1991 -2599
rect -1925 -2565 -1813 -2559
rect -1925 -2599 -1913 -2565
rect -1825 -2599 -1813 -2565
rect -1925 -2605 -1813 -2599
rect -1747 -2565 -1635 -2559
rect -1747 -2599 -1735 -2565
rect -1647 -2599 -1635 -2565
rect -1747 -2605 -1635 -2599
rect -1569 -2565 -1457 -2559
rect -1569 -2599 -1557 -2565
rect -1469 -2599 -1457 -2565
rect -1569 -2605 -1457 -2599
rect -1391 -2565 -1279 -2559
rect -1391 -2599 -1379 -2565
rect -1291 -2599 -1279 -2565
rect -1391 -2605 -1279 -2599
rect -1213 -2565 -1101 -2559
rect -1213 -2599 -1201 -2565
rect -1113 -2599 -1101 -2565
rect -1213 -2605 -1101 -2599
rect -1035 -2565 -923 -2559
rect -1035 -2599 -1023 -2565
rect -935 -2599 -923 -2565
rect -1035 -2605 -923 -2599
rect -857 -2565 -745 -2559
rect -857 -2599 -845 -2565
rect -757 -2599 -745 -2565
rect -857 -2605 -745 -2599
rect -679 -2565 -567 -2559
rect -679 -2599 -667 -2565
rect -579 -2599 -567 -2565
rect -679 -2605 -567 -2599
rect -501 -2565 -389 -2559
rect -501 -2599 -489 -2565
rect -401 -2599 -389 -2565
rect -501 -2605 -389 -2599
rect -323 -2565 -211 -2559
rect -323 -2599 -311 -2565
rect -223 -2599 -211 -2565
rect -323 -2605 -211 -2599
rect -145 -2565 -33 -2559
rect -145 -2599 -133 -2565
rect -45 -2599 -33 -2565
rect -145 -2605 -33 -2599
rect 33 -2565 145 -2559
rect 33 -2599 45 -2565
rect 133 -2599 145 -2565
rect 33 -2605 145 -2599
rect 211 -2565 323 -2559
rect 211 -2599 223 -2565
rect 311 -2599 323 -2565
rect 211 -2605 323 -2599
rect 389 -2565 501 -2559
rect 389 -2599 401 -2565
rect 489 -2599 501 -2565
rect 389 -2605 501 -2599
rect 567 -2565 679 -2559
rect 567 -2599 579 -2565
rect 667 -2599 679 -2565
rect 567 -2605 679 -2599
rect 745 -2565 857 -2559
rect 745 -2599 757 -2565
rect 845 -2599 857 -2565
rect 745 -2605 857 -2599
rect 923 -2565 1035 -2559
rect 923 -2599 935 -2565
rect 1023 -2599 1035 -2565
rect 923 -2605 1035 -2599
rect 1101 -2565 1213 -2559
rect 1101 -2599 1113 -2565
rect 1201 -2599 1213 -2565
rect 1101 -2605 1213 -2599
rect 1279 -2565 1391 -2559
rect 1279 -2599 1291 -2565
rect 1379 -2599 1391 -2565
rect 1279 -2605 1391 -2599
rect 1457 -2565 1569 -2559
rect 1457 -2599 1469 -2565
rect 1557 -2599 1569 -2565
rect 1457 -2605 1569 -2599
rect 1635 -2565 1747 -2559
rect 1635 -2599 1647 -2565
rect 1735 -2599 1747 -2565
rect 1635 -2605 1747 -2599
rect 1813 -2565 1925 -2559
rect 1813 -2599 1825 -2565
rect 1913 -2599 1925 -2565
rect 1813 -2605 1925 -2599
rect 1991 -2565 2103 -2559
rect 1991 -2599 2003 -2565
rect 2091 -2599 2103 -2565
rect 1991 -2605 2103 -2599
rect 2169 -2565 2281 -2559
rect 2169 -2599 2181 -2565
rect 2269 -2599 2281 -2565
rect 2169 -2605 2281 -2599
rect 2347 -2565 2459 -2559
rect 2347 -2599 2359 -2565
rect 2447 -2599 2459 -2565
rect 2347 -2605 2459 -2599
rect 2525 -2565 2637 -2559
rect 2525 -2599 2537 -2565
rect 2625 -2599 2637 -2565
rect 2525 -2605 2637 -2599
rect 2703 -2565 2815 -2559
rect 2703 -2599 2715 -2565
rect 2803 -2599 2815 -2565
rect 2703 -2605 2815 -2599
rect 2881 -2565 2993 -2559
rect 2881 -2599 2893 -2565
rect 2981 -2599 2993 -2565
rect 2881 -2605 2993 -2599
rect 3059 -2565 3171 -2559
rect 3059 -2599 3071 -2565
rect 3159 -2599 3171 -2565
rect 3059 -2605 3171 -2599
rect 3237 -2565 3349 -2559
rect 3237 -2599 3249 -2565
rect 3337 -2599 3349 -2565
rect 3237 -2605 3349 -2599
rect 3415 -2565 3527 -2559
rect 3415 -2599 3427 -2565
rect 3515 -2599 3527 -2565
rect 3415 -2605 3527 -2599
rect 3593 -2565 3705 -2559
rect 3593 -2599 3605 -2565
rect 3693 -2599 3705 -2565
rect 3593 -2605 3705 -2599
rect 3771 -2565 3883 -2559
rect 3771 -2599 3783 -2565
rect 3871 -2599 3883 -2565
rect 3771 -2605 3883 -2599
rect 3949 -2565 4061 -2559
rect 3949 -2599 3961 -2565
rect 4049 -2599 4061 -2565
rect 3949 -2605 4061 -2599
rect 4127 -2565 4239 -2559
rect 4127 -2599 4139 -2565
rect 4227 -2599 4239 -2565
rect 4127 -2605 4239 -2599
rect 4305 -2565 4417 -2559
rect 4305 -2599 4317 -2565
rect 4405 -2599 4417 -2565
rect 4305 -2605 4417 -2599
rect 4483 -2565 4595 -2559
rect 4483 -2599 4495 -2565
rect 4583 -2599 4595 -2565
rect 4483 -2605 4595 -2599
rect 4661 -2565 4773 -2559
rect 4661 -2599 4673 -2565
rect 4761 -2599 4773 -2565
rect 4661 -2605 4773 -2599
rect 4839 -2565 4951 -2559
rect 4839 -2599 4851 -2565
rect 4939 -2599 4951 -2565
rect 4839 -2605 4951 -2599
rect 5017 -2565 5129 -2559
rect 5017 -2599 5029 -2565
rect 5117 -2599 5129 -2565
rect 5017 -2605 5129 -2599
rect 5195 -2565 5307 -2559
rect 5195 -2599 5207 -2565
rect 5295 -2599 5307 -2565
rect 5195 -2605 5307 -2599
rect 5373 -2565 5485 -2559
rect 5373 -2599 5385 -2565
rect 5473 -2599 5485 -2565
rect 5373 -2605 5485 -2599
rect 5551 -2565 5663 -2559
rect 5551 -2599 5563 -2565
rect 5651 -2599 5663 -2565
rect 5551 -2605 5663 -2599
rect 5729 -2565 5841 -2559
rect 5729 -2599 5741 -2565
rect 5829 -2599 5841 -2565
rect 5729 -2605 5841 -2599
rect 5907 -2565 6019 -2559
rect 5907 -2599 5919 -2565
rect 6007 -2599 6019 -2565
rect 5907 -2605 6019 -2599
rect 6085 -2565 6197 -2559
rect 6085 -2599 6097 -2565
rect 6185 -2599 6197 -2565
rect 6085 -2605 6197 -2599
rect 6263 -2565 6375 -2559
rect 6263 -2599 6275 -2565
rect 6363 -2599 6375 -2565
rect 6263 -2605 6375 -2599
rect 6441 -2565 6553 -2559
rect 6441 -2599 6453 -2565
rect 6541 -2599 6553 -2565
rect 6441 -2605 6553 -2599
rect 6619 -2565 6731 -2559
rect 6619 -2599 6631 -2565
rect 6719 -2599 6731 -2565
rect 6619 -2605 6731 -2599
rect 6797 -2565 6909 -2559
rect 6797 -2599 6809 -2565
rect 6897 -2599 6909 -2565
rect 6797 -2605 6909 -2599
rect 6975 -2565 7087 -2559
rect 6975 -2599 6987 -2565
rect 7075 -2599 7087 -2565
rect 6975 -2605 7087 -2599
rect 7153 -2565 7265 -2559
rect 7153 -2599 7165 -2565
rect 7253 -2599 7265 -2565
rect 7153 -2605 7265 -2599
rect 7331 -2565 7443 -2559
rect 7331 -2599 7343 -2565
rect 7431 -2599 7443 -2565
rect 7331 -2605 7443 -2599
rect 7509 -2565 7621 -2559
rect 7509 -2599 7521 -2565
rect 7609 -2599 7621 -2565
rect 7509 -2605 7621 -2599
rect 7687 -2565 7799 -2559
rect 7687 -2599 7699 -2565
rect 7787 -2599 7799 -2565
rect 7687 -2605 7799 -2599
rect 7865 -2565 7977 -2559
rect 7865 -2599 7877 -2565
rect 7965 -2599 7977 -2565
rect 7865 -2605 7977 -2599
rect 8043 -2565 8155 -2559
rect 8043 -2599 8055 -2565
rect 8143 -2599 8155 -2565
rect 8043 -2605 8155 -2599
rect 8221 -2565 8333 -2559
rect 8221 -2599 8233 -2565
rect 8321 -2599 8333 -2565
rect 8221 -2605 8333 -2599
rect 8399 -2565 8511 -2559
rect 8399 -2599 8411 -2565
rect 8499 -2599 8511 -2565
rect 8399 -2605 8511 -2599
rect 8577 -2565 8689 -2559
rect 8577 -2599 8589 -2565
rect 8677 -2599 8689 -2565
rect 8577 -2605 8689 -2599
rect 8755 -2565 8867 -2559
rect 8755 -2599 8767 -2565
rect 8855 -2599 8867 -2565
rect 8755 -2605 8867 -2599
<< properties >>
string FIXED_BBOX -9014 -2684 9014 2684
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 12 l 0.6 m 2 nf 100 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
