magic
tech sky130A
magscale 1 2
timestamp 1723380300
<< error_p >>
rect -5280 1272 -5222 1278
rect -5162 1272 -5104 1278
rect -5044 1272 -4986 1278
rect -4926 1272 -4868 1278
rect -4808 1272 -4750 1278
rect -4690 1272 -4632 1278
rect -4572 1272 -4514 1278
rect -4454 1272 -4396 1278
rect -4336 1272 -4278 1278
rect -4218 1272 -4160 1278
rect -4100 1272 -4042 1278
rect -3982 1272 -3924 1278
rect -3864 1272 -3806 1278
rect -3746 1272 -3688 1278
rect -3628 1272 -3570 1278
rect -3510 1272 -3452 1278
rect -3392 1272 -3334 1278
rect -3274 1272 -3216 1278
rect -3156 1272 -3098 1278
rect -3038 1272 -2980 1278
rect -2920 1272 -2862 1278
rect -2802 1272 -2744 1278
rect -2684 1272 -2626 1278
rect -2566 1272 -2508 1278
rect -2448 1272 -2390 1278
rect -2330 1272 -2272 1278
rect -2212 1272 -2154 1278
rect -2094 1272 -2036 1278
rect -1976 1272 -1918 1278
rect -1858 1272 -1800 1278
rect -1740 1272 -1682 1278
rect -1622 1272 -1564 1278
rect -1504 1272 -1446 1278
rect -1386 1272 -1328 1278
rect -1268 1272 -1210 1278
rect -1150 1272 -1092 1278
rect -1032 1272 -974 1278
rect -914 1272 -856 1278
rect -796 1272 -738 1278
rect -678 1272 -620 1278
rect -560 1272 -502 1278
rect -442 1272 -384 1278
rect -324 1272 -266 1278
rect -206 1272 -148 1278
rect -88 1272 -30 1278
rect 30 1272 88 1278
rect 148 1272 206 1278
rect 266 1272 324 1278
rect 384 1272 442 1278
rect 502 1272 560 1278
rect 620 1272 678 1278
rect 738 1272 796 1278
rect 856 1272 914 1278
rect 974 1272 1032 1278
rect 1092 1272 1150 1278
rect 1210 1272 1268 1278
rect 1328 1272 1386 1278
rect 1446 1272 1504 1278
rect 1564 1272 1622 1278
rect 1682 1272 1740 1278
rect 1800 1272 1858 1278
rect 1918 1272 1976 1278
rect 2036 1272 2094 1278
rect 2154 1272 2212 1278
rect 2272 1272 2330 1278
rect 2390 1272 2448 1278
rect 2508 1272 2566 1278
rect 2626 1272 2684 1278
rect 2744 1272 2802 1278
rect 2862 1272 2920 1278
rect 2980 1272 3038 1278
rect 3098 1272 3156 1278
rect 3216 1272 3274 1278
rect 3334 1272 3392 1278
rect 3452 1272 3510 1278
rect 3570 1272 3628 1278
rect 3688 1272 3746 1278
rect 3806 1272 3864 1278
rect 3924 1272 3982 1278
rect 4042 1272 4100 1278
rect 4160 1272 4218 1278
rect 4278 1272 4336 1278
rect 4396 1272 4454 1278
rect 4514 1272 4572 1278
rect 4632 1272 4690 1278
rect 4750 1272 4808 1278
rect 4868 1272 4926 1278
rect 4986 1272 5044 1278
rect 5104 1272 5162 1278
rect 5222 1272 5280 1278
rect -5280 1238 -5268 1272
rect -5162 1238 -5150 1272
rect -5044 1238 -5032 1272
rect -4926 1238 -4914 1272
rect -4808 1238 -4796 1272
rect -4690 1238 -4678 1272
rect -4572 1238 -4560 1272
rect -4454 1238 -4442 1272
rect -4336 1238 -4324 1272
rect -4218 1238 -4206 1272
rect -4100 1238 -4088 1272
rect -3982 1238 -3970 1272
rect -3864 1238 -3852 1272
rect -3746 1238 -3734 1272
rect -3628 1238 -3616 1272
rect -3510 1238 -3498 1272
rect -3392 1238 -3380 1272
rect -3274 1238 -3262 1272
rect -3156 1238 -3144 1272
rect -3038 1238 -3026 1272
rect -2920 1238 -2908 1272
rect -2802 1238 -2790 1272
rect -2684 1238 -2672 1272
rect -2566 1238 -2554 1272
rect -2448 1238 -2436 1272
rect -2330 1238 -2318 1272
rect -2212 1238 -2200 1272
rect -2094 1238 -2082 1272
rect -1976 1238 -1964 1272
rect -1858 1238 -1846 1272
rect -1740 1238 -1728 1272
rect -1622 1238 -1610 1272
rect -1504 1238 -1492 1272
rect -1386 1238 -1374 1272
rect -1268 1238 -1256 1272
rect -1150 1238 -1138 1272
rect -1032 1238 -1020 1272
rect -914 1238 -902 1272
rect -796 1238 -784 1272
rect -678 1238 -666 1272
rect -560 1238 -548 1272
rect -442 1238 -430 1272
rect -324 1238 -312 1272
rect -206 1238 -194 1272
rect -88 1238 -76 1272
rect 30 1238 42 1272
rect 148 1238 160 1272
rect 266 1238 278 1272
rect 384 1238 396 1272
rect 502 1238 514 1272
rect 620 1238 632 1272
rect 738 1238 750 1272
rect 856 1238 868 1272
rect 974 1238 986 1272
rect 1092 1238 1104 1272
rect 1210 1238 1222 1272
rect 1328 1238 1340 1272
rect 1446 1238 1458 1272
rect 1564 1238 1576 1272
rect 1682 1238 1694 1272
rect 1800 1238 1812 1272
rect 1918 1238 1930 1272
rect 2036 1238 2048 1272
rect 2154 1238 2166 1272
rect 2272 1238 2284 1272
rect 2390 1238 2402 1272
rect 2508 1238 2520 1272
rect 2626 1238 2638 1272
rect 2744 1238 2756 1272
rect 2862 1238 2874 1272
rect 2980 1238 2992 1272
rect 3098 1238 3110 1272
rect 3216 1238 3228 1272
rect 3334 1238 3346 1272
rect 3452 1238 3464 1272
rect 3570 1238 3582 1272
rect 3688 1238 3700 1272
rect 3806 1238 3818 1272
rect 3924 1238 3936 1272
rect 4042 1238 4054 1272
rect 4160 1238 4172 1272
rect 4278 1238 4290 1272
rect 4396 1238 4408 1272
rect 4514 1238 4526 1272
rect 4632 1238 4644 1272
rect 4750 1238 4762 1272
rect 4868 1238 4880 1272
rect 4986 1238 4998 1272
rect 5104 1238 5116 1272
rect 5222 1238 5234 1272
rect -5280 1232 -5222 1238
rect -5162 1232 -5104 1238
rect -5044 1232 -4986 1238
rect -4926 1232 -4868 1238
rect -4808 1232 -4750 1238
rect -4690 1232 -4632 1238
rect -4572 1232 -4514 1238
rect -4454 1232 -4396 1238
rect -4336 1232 -4278 1238
rect -4218 1232 -4160 1238
rect -4100 1232 -4042 1238
rect -3982 1232 -3924 1238
rect -3864 1232 -3806 1238
rect -3746 1232 -3688 1238
rect -3628 1232 -3570 1238
rect -3510 1232 -3452 1238
rect -3392 1232 -3334 1238
rect -3274 1232 -3216 1238
rect -3156 1232 -3098 1238
rect -3038 1232 -2980 1238
rect -2920 1232 -2862 1238
rect -2802 1232 -2744 1238
rect -2684 1232 -2626 1238
rect -2566 1232 -2508 1238
rect -2448 1232 -2390 1238
rect -2330 1232 -2272 1238
rect -2212 1232 -2154 1238
rect -2094 1232 -2036 1238
rect -1976 1232 -1918 1238
rect -1858 1232 -1800 1238
rect -1740 1232 -1682 1238
rect -1622 1232 -1564 1238
rect -1504 1232 -1446 1238
rect -1386 1232 -1328 1238
rect -1268 1232 -1210 1238
rect -1150 1232 -1092 1238
rect -1032 1232 -974 1238
rect -914 1232 -856 1238
rect -796 1232 -738 1238
rect -678 1232 -620 1238
rect -560 1232 -502 1238
rect -442 1232 -384 1238
rect -324 1232 -266 1238
rect -206 1232 -148 1238
rect -88 1232 -30 1238
rect 30 1232 88 1238
rect 148 1232 206 1238
rect 266 1232 324 1238
rect 384 1232 442 1238
rect 502 1232 560 1238
rect 620 1232 678 1238
rect 738 1232 796 1238
rect 856 1232 914 1238
rect 974 1232 1032 1238
rect 1092 1232 1150 1238
rect 1210 1232 1268 1238
rect 1328 1232 1386 1238
rect 1446 1232 1504 1238
rect 1564 1232 1622 1238
rect 1682 1232 1740 1238
rect 1800 1232 1858 1238
rect 1918 1232 1976 1238
rect 2036 1232 2094 1238
rect 2154 1232 2212 1238
rect 2272 1232 2330 1238
rect 2390 1232 2448 1238
rect 2508 1232 2566 1238
rect 2626 1232 2684 1238
rect 2744 1232 2802 1238
rect 2862 1232 2920 1238
rect 2980 1232 3038 1238
rect 3098 1232 3156 1238
rect 3216 1232 3274 1238
rect 3334 1232 3392 1238
rect 3452 1232 3510 1238
rect 3570 1232 3628 1238
rect 3688 1232 3746 1238
rect 3806 1232 3864 1238
rect 3924 1232 3982 1238
rect 4042 1232 4100 1238
rect 4160 1232 4218 1238
rect 4278 1232 4336 1238
rect 4396 1232 4454 1238
rect 4514 1232 4572 1238
rect 4632 1232 4690 1238
rect 4750 1232 4808 1238
rect 4868 1232 4926 1238
rect 4986 1232 5044 1238
rect 5104 1232 5162 1238
rect 5222 1232 5280 1238
rect -5280 -1238 -5222 -1232
rect -5162 -1238 -5104 -1232
rect -5044 -1238 -4986 -1232
rect -4926 -1238 -4868 -1232
rect -4808 -1238 -4750 -1232
rect -4690 -1238 -4632 -1232
rect -4572 -1238 -4514 -1232
rect -4454 -1238 -4396 -1232
rect -4336 -1238 -4278 -1232
rect -4218 -1238 -4160 -1232
rect -4100 -1238 -4042 -1232
rect -3982 -1238 -3924 -1232
rect -3864 -1238 -3806 -1232
rect -3746 -1238 -3688 -1232
rect -3628 -1238 -3570 -1232
rect -3510 -1238 -3452 -1232
rect -3392 -1238 -3334 -1232
rect -3274 -1238 -3216 -1232
rect -3156 -1238 -3098 -1232
rect -3038 -1238 -2980 -1232
rect -2920 -1238 -2862 -1232
rect -2802 -1238 -2744 -1232
rect -2684 -1238 -2626 -1232
rect -2566 -1238 -2508 -1232
rect -2448 -1238 -2390 -1232
rect -2330 -1238 -2272 -1232
rect -2212 -1238 -2154 -1232
rect -2094 -1238 -2036 -1232
rect -1976 -1238 -1918 -1232
rect -1858 -1238 -1800 -1232
rect -1740 -1238 -1682 -1232
rect -1622 -1238 -1564 -1232
rect -1504 -1238 -1446 -1232
rect -1386 -1238 -1328 -1232
rect -1268 -1238 -1210 -1232
rect -1150 -1238 -1092 -1232
rect -1032 -1238 -974 -1232
rect -914 -1238 -856 -1232
rect -796 -1238 -738 -1232
rect -678 -1238 -620 -1232
rect -560 -1238 -502 -1232
rect -442 -1238 -384 -1232
rect -324 -1238 -266 -1232
rect -206 -1238 -148 -1232
rect -88 -1238 -30 -1232
rect 30 -1238 88 -1232
rect 148 -1238 206 -1232
rect 266 -1238 324 -1232
rect 384 -1238 442 -1232
rect 502 -1238 560 -1232
rect 620 -1238 678 -1232
rect 738 -1238 796 -1232
rect 856 -1238 914 -1232
rect 974 -1238 1032 -1232
rect 1092 -1238 1150 -1232
rect 1210 -1238 1268 -1232
rect 1328 -1238 1386 -1232
rect 1446 -1238 1504 -1232
rect 1564 -1238 1622 -1232
rect 1682 -1238 1740 -1232
rect 1800 -1238 1858 -1232
rect 1918 -1238 1976 -1232
rect 2036 -1238 2094 -1232
rect 2154 -1238 2212 -1232
rect 2272 -1238 2330 -1232
rect 2390 -1238 2448 -1232
rect 2508 -1238 2566 -1232
rect 2626 -1238 2684 -1232
rect 2744 -1238 2802 -1232
rect 2862 -1238 2920 -1232
rect 2980 -1238 3038 -1232
rect 3098 -1238 3156 -1232
rect 3216 -1238 3274 -1232
rect 3334 -1238 3392 -1232
rect 3452 -1238 3510 -1232
rect 3570 -1238 3628 -1232
rect 3688 -1238 3746 -1232
rect 3806 -1238 3864 -1232
rect 3924 -1238 3982 -1232
rect 4042 -1238 4100 -1232
rect 4160 -1238 4218 -1232
rect 4278 -1238 4336 -1232
rect 4396 -1238 4454 -1232
rect 4514 -1238 4572 -1232
rect 4632 -1238 4690 -1232
rect 4750 -1238 4808 -1232
rect 4868 -1238 4926 -1232
rect 4986 -1238 5044 -1232
rect 5104 -1238 5162 -1232
rect 5222 -1238 5280 -1232
rect -5280 -1272 -5268 -1238
rect -5162 -1272 -5150 -1238
rect -5044 -1272 -5032 -1238
rect -4926 -1272 -4914 -1238
rect -4808 -1272 -4796 -1238
rect -4690 -1272 -4678 -1238
rect -4572 -1272 -4560 -1238
rect -4454 -1272 -4442 -1238
rect -4336 -1272 -4324 -1238
rect -4218 -1272 -4206 -1238
rect -4100 -1272 -4088 -1238
rect -3982 -1272 -3970 -1238
rect -3864 -1272 -3852 -1238
rect -3746 -1272 -3734 -1238
rect -3628 -1272 -3616 -1238
rect -3510 -1272 -3498 -1238
rect -3392 -1272 -3380 -1238
rect -3274 -1272 -3262 -1238
rect -3156 -1272 -3144 -1238
rect -3038 -1272 -3026 -1238
rect -2920 -1272 -2908 -1238
rect -2802 -1272 -2790 -1238
rect -2684 -1272 -2672 -1238
rect -2566 -1272 -2554 -1238
rect -2448 -1272 -2436 -1238
rect -2330 -1272 -2318 -1238
rect -2212 -1272 -2200 -1238
rect -2094 -1272 -2082 -1238
rect -1976 -1272 -1964 -1238
rect -1858 -1272 -1846 -1238
rect -1740 -1272 -1728 -1238
rect -1622 -1272 -1610 -1238
rect -1504 -1272 -1492 -1238
rect -1386 -1272 -1374 -1238
rect -1268 -1272 -1256 -1238
rect -1150 -1272 -1138 -1238
rect -1032 -1272 -1020 -1238
rect -914 -1272 -902 -1238
rect -796 -1272 -784 -1238
rect -678 -1272 -666 -1238
rect -560 -1272 -548 -1238
rect -442 -1272 -430 -1238
rect -324 -1272 -312 -1238
rect -206 -1272 -194 -1238
rect -88 -1272 -76 -1238
rect 30 -1272 42 -1238
rect 148 -1272 160 -1238
rect 266 -1272 278 -1238
rect 384 -1272 396 -1238
rect 502 -1272 514 -1238
rect 620 -1272 632 -1238
rect 738 -1272 750 -1238
rect 856 -1272 868 -1238
rect 974 -1272 986 -1238
rect 1092 -1272 1104 -1238
rect 1210 -1272 1222 -1238
rect 1328 -1272 1340 -1238
rect 1446 -1272 1458 -1238
rect 1564 -1272 1576 -1238
rect 1682 -1272 1694 -1238
rect 1800 -1272 1812 -1238
rect 1918 -1272 1930 -1238
rect 2036 -1272 2048 -1238
rect 2154 -1272 2166 -1238
rect 2272 -1272 2284 -1238
rect 2390 -1272 2402 -1238
rect 2508 -1272 2520 -1238
rect 2626 -1272 2638 -1238
rect 2744 -1272 2756 -1238
rect 2862 -1272 2874 -1238
rect 2980 -1272 2992 -1238
rect 3098 -1272 3110 -1238
rect 3216 -1272 3228 -1238
rect 3334 -1272 3346 -1238
rect 3452 -1272 3464 -1238
rect 3570 -1272 3582 -1238
rect 3688 -1272 3700 -1238
rect 3806 -1272 3818 -1238
rect 3924 -1272 3936 -1238
rect 4042 -1272 4054 -1238
rect 4160 -1272 4172 -1238
rect 4278 -1272 4290 -1238
rect 4396 -1272 4408 -1238
rect 4514 -1272 4526 -1238
rect 4632 -1272 4644 -1238
rect 4750 -1272 4762 -1238
rect 4868 -1272 4880 -1238
rect 4986 -1272 4998 -1238
rect 5104 -1272 5116 -1238
rect 5222 -1272 5234 -1238
rect -5280 -1278 -5222 -1272
rect -5162 -1278 -5104 -1272
rect -5044 -1278 -4986 -1272
rect -4926 -1278 -4868 -1272
rect -4808 -1278 -4750 -1272
rect -4690 -1278 -4632 -1272
rect -4572 -1278 -4514 -1272
rect -4454 -1278 -4396 -1272
rect -4336 -1278 -4278 -1272
rect -4218 -1278 -4160 -1272
rect -4100 -1278 -4042 -1272
rect -3982 -1278 -3924 -1272
rect -3864 -1278 -3806 -1272
rect -3746 -1278 -3688 -1272
rect -3628 -1278 -3570 -1272
rect -3510 -1278 -3452 -1272
rect -3392 -1278 -3334 -1272
rect -3274 -1278 -3216 -1272
rect -3156 -1278 -3098 -1272
rect -3038 -1278 -2980 -1272
rect -2920 -1278 -2862 -1272
rect -2802 -1278 -2744 -1272
rect -2684 -1278 -2626 -1272
rect -2566 -1278 -2508 -1272
rect -2448 -1278 -2390 -1272
rect -2330 -1278 -2272 -1272
rect -2212 -1278 -2154 -1272
rect -2094 -1278 -2036 -1272
rect -1976 -1278 -1918 -1272
rect -1858 -1278 -1800 -1272
rect -1740 -1278 -1682 -1272
rect -1622 -1278 -1564 -1272
rect -1504 -1278 -1446 -1272
rect -1386 -1278 -1328 -1272
rect -1268 -1278 -1210 -1272
rect -1150 -1278 -1092 -1272
rect -1032 -1278 -974 -1272
rect -914 -1278 -856 -1272
rect -796 -1278 -738 -1272
rect -678 -1278 -620 -1272
rect -560 -1278 -502 -1272
rect -442 -1278 -384 -1272
rect -324 -1278 -266 -1272
rect -206 -1278 -148 -1272
rect -88 -1278 -30 -1272
rect 30 -1278 88 -1272
rect 148 -1278 206 -1272
rect 266 -1278 324 -1272
rect 384 -1278 442 -1272
rect 502 -1278 560 -1272
rect 620 -1278 678 -1272
rect 738 -1278 796 -1272
rect 856 -1278 914 -1272
rect 974 -1278 1032 -1272
rect 1092 -1278 1150 -1272
rect 1210 -1278 1268 -1272
rect 1328 -1278 1386 -1272
rect 1446 -1278 1504 -1272
rect 1564 -1278 1622 -1272
rect 1682 -1278 1740 -1272
rect 1800 -1278 1858 -1272
rect 1918 -1278 1976 -1272
rect 2036 -1278 2094 -1272
rect 2154 -1278 2212 -1272
rect 2272 -1278 2330 -1272
rect 2390 -1278 2448 -1272
rect 2508 -1278 2566 -1272
rect 2626 -1278 2684 -1272
rect 2744 -1278 2802 -1272
rect 2862 -1278 2920 -1272
rect 2980 -1278 3038 -1272
rect 3098 -1278 3156 -1272
rect 3216 -1278 3274 -1272
rect 3334 -1278 3392 -1272
rect 3452 -1278 3510 -1272
rect 3570 -1278 3628 -1272
rect 3688 -1278 3746 -1272
rect 3806 -1278 3864 -1272
rect 3924 -1278 3982 -1272
rect 4042 -1278 4100 -1272
rect 4160 -1278 4218 -1272
rect 4278 -1278 4336 -1272
rect 4396 -1278 4454 -1272
rect 4514 -1278 4572 -1272
rect 4632 -1278 4690 -1272
rect 4750 -1278 4808 -1272
rect 4868 -1278 4926 -1272
rect 4986 -1278 5044 -1272
rect 5104 -1278 5162 -1272
rect 5222 -1278 5280 -1272
<< pwell >>
rect -5477 -1410 5477 1410
<< nmos >>
rect -5281 -1200 -5221 1200
rect -5163 -1200 -5103 1200
rect -5045 -1200 -4985 1200
rect -4927 -1200 -4867 1200
rect -4809 -1200 -4749 1200
rect -4691 -1200 -4631 1200
rect -4573 -1200 -4513 1200
rect -4455 -1200 -4395 1200
rect -4337 -1200 -4277 1200
rect -4219 -1200 -4159 1200
rect -4101 -1200 -4041 1200
rect -3983 -1200 -3923 1200
rect -3865 -1200 -3805 1200
rect -3747 -1200 -3687 1200
rect -3629 -1200 -3569 1200
rect -3511 -1200 -3451 1200
rect -3393 -1200 -3333 1200
rect -3275 -1200 -3215 1200
rect -3157 -1200 -3097 1200
rect -3039 -1200 -2979 1200
rect -2921 -1200 -2861 1200
rect -2803 -1200 -2743 1200
rect -2685 -1200 -2625 1200
rect -2567 -1200 -2507 1200
rect -2449 -1200 -2389 1200
rect -2331 -1200 -2271 1200
rect -2213 -1200 -2153 1200
rect -2095 -1200 -2035 1200
rect -1977 -1200 -1917 1200
rect -1859 -1200 -1799 1200
rect -1741 -1200 -1681 1200
rect -1623 -1200 -1563 1200
rect -1505 -1200 -1445 1200
rect -1387 -1200 -1327 1200
rect -1269 -1200 -1209 1200
rect -1151 -1200 -1091 1200
rect -1033 -1200 -973 1200
rect -915 -1200 -855 1200
rect -797 -1200 -737 1200
rect -679 -1200 -619 1200
rect -561 -1200 -501 1200
rect -443 -1200 -383 1200
rect -325 -1200 -265 1200
rect -207 -1200 -147 1200
rect -89 -1200 -29 1200
rect 29 -1200 89 1200
rect 147 -1200 207 1200
rect 265 -1200 325 1200
rect 383 -1200 443 1200
rect 501 -1200 561 1200
rect 619 -1200 679 1200
rect 737 -1200 797 1200
rect 855 -1200 915 1200
rect 973 -1200 1033 1200
rect 1091 -1200 1151 1200
rect 1209 -1200 1269 1200
rect 1327 -1200 1387 1200
rect 1445 -1200 1505 1200
rect 1563 -1200 1623 1200
rect 1681 -1200 1741 1200
rect 1799 -1200 1859 1200
rect 1917 -1200 1977 1200
rect 2035 -1200 2095 1200
rect 2153 -1200 2213 1200
rect 2271 -1200 2331 1200
rect 2389 -1200 2449 1200
rect 2507 -1200 2567 1200
rect 2625 -1200 2685 1200
rect 2743 -1200 2803 1200
rect 2861 -1200 2921 1200
rect 2979 -1200 3039 1200
rect 3097 -1200 3157 1200
rect 3215 -1200 3275 1200
rect 3333 -1200 3393 1200
rect 3451 -1200 3511 1200
rect 3569 -1200 3629 1200
rect 3687 -1200 3747 1200
rect 3805 -1200 3865 1200
rect 3923 -1200 3983 1200
rect 4041 -1200 4101 1200
rect 4159 -1200 4219 1200
rect 4277 -1200 4337 1200
rect 4395 -1200 4455 1200
rect 4513 -1200 4573 1200
rect 4631 -1200 4691 1200
rect 4749 -1200 4809 1200
rect 4867 -1200 4927 1200
rect 4985 -1200 5045 1200
rect 5103 -1200 5163 1200
rect 5221 -1200 5281 1200
<< ndiff >>
rect -5339 1188 -5281 1200
rect -5339 -1188 -5327 1188
rect -5293 -1188 -5281 1188
rect -5339 -1200 -5281 -1188
rect -5221 1188 -5163 1200
rect -5221 -1188 -5209 1188
rect -5175 -1188 -5163 1188
rect -5221 -1200 -5163 -1188
rect -5103 1188 -5045 1200
rect -5103 -1188 -5091 1188
rect -5057 -1188 -5045 1188
rect -5103 -1200 -5045 -1188
rect -4985 1188 -4927 1200
rect -4985 -1188 -4973 1188
rect -4939 -1188 -4927 1188
rect -4985 -1200 -4927 -1188
rect -4867 1188 -4809 1200
rect -4867 -1188 -4855 1188
rect -4821 -1188 -4809 1188
rect -4867 -1200 -4809 -1188
rect -4749 1188 -4691 1200
rect -4749 -1188 -4737 1188
rect -4703 -1188 -4691 1188
rect -4749 -1200 -4691 -1188
rect -4631 1188 -4573 1200
rect -4631 -1188 -4619 1188
rect -4585 -1188 -4573 1188
rect -4631 -1200 -4573 -1188
rect -4513 1188 -4455 1200
rect -4513 -1188 -4501 1188
rect -4467 -1188 -4455 1188
rect -4513 -1200 -4455 -1188
rect -4395 1188 -4337 1200
rect -4395 -1188 -4383 1188
rect -4349 -1188 -4337 1188
rect -4395 -1200 -4337 -1188
rect -4277 1188 -4219 1200
rect -4277 -1188 -4265 1188
rect -4231 -1188 -4219 1188
rect -4277 -1200 -4219 -1188
rect -4159 1188 -4101 1200
rect -4159 -1188 -4147 1188
rect -4113 -1188 -4101 1188
rect -4159 -1200 -4101 -1188
rect -4041 1188 -3983 1200
rect -4041 -1188 -4029 1188
rect -3995 -1188 -3983 1188
rect -4041 -1200 -3983 -1188
rect -3923 1188 -3865 1200
rect -3923 -1188 -3911 1188
rect -3877 -1188 -3865 1188
rect -3923 -1200 -3865 -1188
rect -3805 1188 -3747 1200
rect -3805 -1188 -3793 1188
rect -3759 -1188 -3747 1188
rect -3805 -1200 -3747 -1188
rect -3687 1188 -3629 1200
rect -3687 -1188 -3675 1188
rect -3641 -1188 -3629 1188
rect -3687 -1200 -3629 -1188
rect -3569 1188 -3511 1200
rect -3569 -1188 -3557 1188
rect -3523 -1188 -3511 1188
rect -3569 -1200 -3511 -1188
rect -3451 1188 -3393 1200
rect -3451 -1188 -3439 1188
rect -3405 -1188 -3393 1188
rect -3451 -1200 -3393 -1188
rect -3333 1188 -3275 1200
rect -3333 -1188 -3321 1188
rect -3287 -1188 -3275 1188
rect -3333 -1200 -3275 -1188
rect -3215 1188 -3157 1200
rect -3215 -1188 -3203 1188
rect -3169 -1188 -3157 1188
rect -3215 -1200 -3157 -1188
rect -3097 1188 -3039 1200
rect -3097 -1188 -3085 1188
rect -3051 -1188 -3039 1188
rect -3097 -1200 -3039 -1188
rect -2979 1188 -2921 1200
rect -2979 -1188 -2967 1188
rect -2933 -1188 -2921 1188
rect -2979 -1200 -2921 -1188
rect -2861 1188 -2803 1200
rect -2861 -1188 -2849 1188
rect -2815 -1188 -2803 1188
rect -2861 -1200 -2803 -1188
rect -2743 1188 -2685 1200
rect -2743 -1188 -2731 1188
rect -2697 -1188 -2685 1188
rect -2743 -1200 -2685 -1188
rect -2625 1188 -2567 1200
rect -2625 -1188 -2613 1188
rect -2579 -1188 -2567 1188
rect -2625 -1200 -2567 -1188
rect -2507 1188 -2449 1200
rect -2507 -1188 -2495 1188
rect -2461 -1188 -2449 1188
rect -2507 -1200 -2449 -1188
rect -2389 1188 -2331 1200
rect -2389 -1188 -2377 1188
rect -2343 -1188 -2331 1188
rect -2389 -1200 -2331 -1188
rect -2271 1188 -2213 1200
rect -2271 -1188 -2259 1188
rect -2225 -1188 -2213 1188
rect -2271 -1200 -2213 -1188
rect -2153 1188 -2095 1200
rect -2153 -1188 -2141 1188
rect -2107 -1188 -2095 1188
rect -2153 -1200 -2095 -1188
rect -2035 1188 -1977 1200
rect -2035 -1188 -2023 1188
rect -1989 -1188 -1977 1188
rect -2035 -1200 -1977 -1188
rect -1917 1188 -1859 1200
rect -1917 -1188 -1905 1188
rect -1871 -1188 -1859 1188
rect -1917 -1200 -1859 -1188
rect -1799 1188 -1741 1200
rect -1799 -1188 -1787 1188
rect -1753 -1188 -1741 1188
rect -1799 -1200 -1741 -1188
rect -1681 1188 -1623 1200
rect -1681 -1188 -1669 1188
rect -1635 -1188 -1623 1188
rect -1681 -1200 -1623 -1188
rect -1563 1188 -1505 1200
rect -1563 -1188 -1551 1188
rect -1517 -1188 -1505 1188
rect -1563 -1200 -1505 -1188
rect -1445 1188 -1387 1200
rect -1445 -1188 -1433 1188
rect -1399 -1188 -1387 1188
rect -1445 -1200 -1387 -1188
rect -1327 1188 -1269 1200
rect -1327 -1188 -1315 1188
rect -1281 -1188 -1269 1188
rect -1327 -1200 -1269 -1188
rect -1209 1188 -1151 1200
rect -1209 -1188 -1197 1188
rect -1163 -1188 -1151 1188
rect -1209 -1200 -1151 -1188
rect -1091 1188 -1033 1200
rect -1091 -1188 -1079 1188
rect -1045 -1188 -1033 1188
rect -1091 -1200 -1033 -1188
rect -973 1188 -915 1200
rect -973 -1188 -961 1188
rect -927 -1188 -915 1188
rect -973 -1200 -915 -1188
rect -855 1188 -797 1200
rect -855 -1188 -843 1188
rect -809 -1188 -797 1188
rect -855 -1200 -797 -1188
rect -737 1188 -679 1200
rect -737 -1188 -725 1188
rect -691 -1188 -679 1188
rect -737 -1200 -679 -1188
rect -619 1188 -561 1200
rect -619 -1188 -607 1188
rect -573 -1188 -561 1188
rect -619 -1200 -561 -1188
rect -501 1188 -443 1200
rect -501 -1188 -489 1188
rect -455 -1188 -443 1188
rect -501 -1200 -443 -1188
rect -383 1188 -325 1200
rect -383 -1188 -371 1188
rect -337 -1188 -325 1188
rect -383 -1200 -325 -1188
rect -265 1188 -207 1200
rect -265 -1188 -253 1188
rect -219 -1188 -207 1188
rect -265 -1200 -207 -1188
rect -147 1188 -89 1200
rect -147 -1188 -135 1188
rect -101 -1188 -89 1188
rect -147 -1200 -89 -1188
rect -29 1188 29 1200
rect -29 -1188 -17 1188
rect 17 -1188 29 1188
rect -29 -1200 29 -1188
rect 89 1188 147 1200
rect 89 -1188 101 1188
rect 135 -1188 147 1188
rect 89 -1200 147 -1188
rect 207 1188 265 1200
rect 207 -1188 219 1188
rect 253 -1188 265 1188
rect 207 -1200 265 -1188
rect 325 1188 383 1200
rect 325 -1188 337 1188
rect 371 -1188 383 1188
rect 325 -1200 383 -1188
rect 443 1188 501 1200
rect 443 -1188 455 1188
rect 489 -1188 501 1188
rect 443 -1200 501 -1188
rect 561 1188 619 1200
rect 561 -1188 573 1188
rect 607 -1188 619 1188
rect 561 -1200 619 -1188
rect 679 1188 737 1200
rect 679 -1188 691 1188
rect 725 -1188 737 1188
rect 679 -1200 737 -1188
rect 797 1188 855 1200
rect 797 -1188 809 1188
rect 843 -1188 855 1188
rect 797 -1200 855 -1188
rect 915 1188 973 1200
rect 915 -1188 927 1188
rect 961 -1188 973 1188
rect 915 -1200 973 -1188
rect 1033 1188 1091 1200
rect 1033 -1188 1045 1188
rect 1079 -1188 1091 1188
rect 1033 -1200 1091 -1188
rect 1151 1188 1209 1200
rect 1151 -1188 1163 1188
rect 1197 -1188 1209 1188
rect 1151 -1200 1209 -1188
rect 1269 1188 1327 1200
rect 1269 -1188 1281 1188
rect 1315 -1188 1327 1188
rect 1269 -1200 1327 -1188
rect 1387 1188 1445 1200
rect 1387 -1188 1399 1188
rect 1433 -1188 1445 1188
rect 1387 -1200 1445 -1188
rect 1505 1188 1563 1200
rect 1505 -1188 1517 1188
rect 1551 -1188 1563 1188
rect 1505 -1200 1563 -1188
rect 1623 1188 1681 1200
rect 1623 -1188 1635 1188
rect 1669 -1188 1681 1188
rect 1623 -1200 1681 -1188
rect 1741 1188 1799 1200
rect 1741 -1188 1753 1188
rect 1787 -1188 1799 1188
rect 1741 -1200 1799 -1188
rect 1859 1188 1917 1200
rect 1859 -1188 1871 1188
rect 1905 -1188 1917 1188
rect 1859 -1200 1917 -1188
rect 1977 1188 2035 1200
rect 1977 -1188 1989 1188
rect 2023 -1188 2035 1188
rect 1977 -1200 2035 -1188
rect 2095 1188 2153 1200
rect 2095 -1188 2107 1188
rect 2141 -1188 2153 1188
rect 2095 -1200 2153 -1188
rect 2213 1188 2271 1200
rect 2213 -1188 2225 1188
rect 2259 -1188 2271 1188
rect 2213 -1200 2271 -1188
rect 2331 1188 2389 1200
rect 2331 -1188 2343 1188
rect 2377 -1188 2389 1188
rect 2331 -1200 2389 -1188
rect 2449 1188 2507 1200
rect 2449 -1188 2461 1188
rect 2495 -1188 2507 1188
rect 2449 -1200 2507 -1188
rect 2567 1188 2625 1200
rect 2567 -1188 2579 1188
rect 2613 -1188 2625 1188
rect 2567 -1200 2625 -1188
rect 2685 1188 2743 1200
rect 2685 -1188 2697 1188
rect 2731 -1188 2743 1188
rect 2685 -1200 2743 -1188
rect 2803 1188 2861 1200
rect 2803 -1188 2815 1188
rect 2849 -1188 2861 1188
rect 2803 -1200 2861 -1188
rect 2921 1188 2979 1200
rect 2921 -1188 2933 1188
rect 2967 -1188 2979 1188
rect 2921 -1200 2979 -1188
rect 3039 1188 3097 1200
rect 3039 -1188 3051 1188
rect 3085 -1188 3097 1188
rect 3039 -1200 3097 -1188
rect 3157 1188 3215 1200
rect 3157 -1188 3169 1188
rect 3203 -1188 3215 1188
rect 3157 -1200 3215 -1188
rect 3275 1188 3333 1200
rect 3275 -1188 3287 1188
rect 3321 -1188 3333 1188
rect 3275 -1200 3333 -1188
rect 3393 1188 3451 1200
rect 3393 -1188 3405 1188
rect 3439 -1188 3451 1188
rect 3393 -1200 3451 -1188
rect 3511 1188 3569 1200
rect 3511 -1188 3523 1188
rect 3557 -1188 3569 1188
rect 3511 -1200 3569 -1188
rect 3629 1188 3687 1200
rect 3629 -1188 3641 1188
rect 3675 -1188 3687 1188
rect 3629 -1200 3687 -1188
rect 3747 1188 3805 1200
rect 3747 -1188 3759 1188
rect 3793 -1188 3805 1188
rect 3747 -1200 3805 -1188
rect 3865 1188 3923 1200
rect 3865 -1188 3877 1188
rect 3911 -1188 3923 1188
rect 3865 -1200 3923 -1188
rect 3983 1188 4041 1200
rect 3983 -1188 3995 1188
rect 4029 -1188 4041 1188
rect 3983 -1200 4041 -1188
rect 4101 1188 4159 1200
rect 4101 -1188 4113 1188
rect 4147 -1188 4159 1188
rect 4101 -1200 4159 -1188
rect 4219 1188 4277 1200
rect 4219 -1188 4231 1188
rect 4265 -1188 4277 1188
rect 4219 -1200 4277 -1188
rect 4337 1188 4395 1200
rect 4337 -1188 4349 1188
rect 4383 -1188 4395 1188
rect 4337 -1200 4395 -1188
rect 4455 1188 4513 1200
rect 4455 -1188 4467 1188
rect 4501 -1188 4513 1188
rect 4455 -1200 4513 -1188
rect 4573 1188 4631 1200
rect 4573 -1188 4585 1188
rect 4619 -1188 4631 1188
rect 4573 -1200 4631 -1188
rect 4691 1188 4749 1200
rect 4691 -1188 4703 1188
rect 4737 -1188 4749 1188
rect 4691 -1200 4749 -1188
rect 4809 1188 4867 1200
rect 4809 -1188 4821 1188
rect 4855 -1188 4867 1188
rect 4809 -1200 4867 -1188
rect 4927 1188 4985 1200
rect 4927 -1188 4939 1188
rect 4973 -1188 4985 1188
rect 4927 -1200 4985 -1188
rect 5045 1188 5103 1200
rect 5045 -1188 5057 1188
rect 5091 -1188 5103 1188
rect 5045 -1200 5103 -1188
rect 5163 1188 5221 1200
rect 5163 -1188 5175 1188
rect 5209 -1188 5221 1188
rect 5163 -1200 5221 -1188
rect 5281 1188 5339 1200
rect 5281 -1188 5293 1188
rect 5327 -1188 5339 1188
rect 5281 -1200 5339 -1188
<< ndiffc >>
rect -5327 -1188 -5293 1188
rect -5209 -1188 -5175 1188
rect -5091 -1188 -5057 1188
rect -4973 -1188 -4939 1188
rect -4855 -1188 -4821 1188
rect -4737 -1188 -4703 1188
rect -4619 -1188 -4585 1188
rect -4501 -1188 -4467 1188
rect -4383 -1188 -4349 1188
rect -4265 -1188 -4231 1188
rect -4147 -1188 -4113 1188
rect -4029 -1188 -3995 1188
rect -3911 -1188 -3877 1188
rect -3793 -1188 -3759 1188
rect -3675 -1188 -3641 1188
rect -3557 -1188 -3523 1188
rect -3439 -1188 -3405 1188
rect -3321 -1188 -3287 1188
rect -3203 -1188 -3169 1188
rect -3085 -1188 -3051 1188
rect -2967 -1188 -2933 1188
rect -2849 -1188 -2815 1188
rect -2731 -1188 -2697 1188
rect -2613 -1188 -2579 1188
rect -2495 -1188 -2461 1188
rect -2377 -1188 -2343 1188
rect -2259 -1188 -2225 1188
rect -2141 -1188 -2107 1188
rect -2023 -1188 -1989 1188
rect -1905 -1188 -1871 1188
rect -1787 -1188 -1753 1188
rect -1669 -1188 -1635 1188
rect -1551 -1188 -1517 1188
rect -1433 -1188 -1399 1188
rect -1315 -1188 -1281 1188
rect -1197 -1188 -1163 1188
rect -1079 -1188 -1045 1188
rect -961 -1188 -927 1188
rect -843 -1188 -809 1188
rect -725 -1188 -691 1188
rect -607 -1188 -573 1188
rect -489 -1188 -455 1188
rect -371 -1188 -337 1188
rect -253 -1188 -219 1188
rect -135 -1188 -101 1188
rect -17 -1188 17 1188
rect 101 -1188 135 1188
rect 219 -1188 253 1188
rect 337 -1188 371 1188
rect 455 -1188 489 1188
rect 573 -1188 607 1188
rect 691 -1188 725 1188
rect 809 -1188 843 1188
rect 927 -1188 961 1188
rect 1045 -1188 1079 1188
rect 1163 -1188 1197 1188
rect 1281 -1188 1315 1188
rect 1399 -1188 1433 1188
rect 1517 -1188 1551 1188
rect 1635 -1188 1669 1188
rect 1753 -1188 1787 1188
rect 1871 -1188 1905 1188
rect 1989 -1188 2023 1188
rect 2107 -1188 2141 1188
rect 2225 -1188 2259 1188
rect 2343 -1188 2377 1188
rect 2461 -1188 2495 1188
rect 2579 -1188 2613 1188
rect 2697 -1188 2731 1188
rect 2815 -1188 2849 1188
rect 2933 -1188 2967 1188
rect 3051 -1188 3085 1188
rect 3169 -1188 3203 1188
rect 3287 -1188 3321 1188
rect 3405 -1188 3439 1188
rect 3523 -1188 3557 1188
rect 3641 -1188 3675 1188
rect 3759 -1188 3793 1188
rect 3877 -1188 3911 1188
rect 3995 -1188 4029 1188
rect 4113 -1188 4147 1188
rect 4231 -1188 4265 1188
rect 4349 -1188 4383 1188
rect 4467 -1188 4501 1188
rect 4585 -1188 4619 1188
rect 4703 -1188 4737 1188
rect 4821 -1188 4855 1188
rect 4939 -1188 4973 1188
rect 5057 -1188 5091 1188
rect 5175 -1188 5209 1188
rect 5293 -1188 5327 1188
<< psubdiff >>
rect -5441 1340 -5345 1374
rect 5345 1340 5441 1374
rect -5441 1278 -5407 1340
rect 5407 1278 5441 1340
rect -5441 -1340 -5407 -1278
rect 5407 -1340 5441 -1278
rect -5441 -1374 -5345 -1340
rect 5345 -1374 5441 -1340
<< psubdiffcont >>
rect -5345 1340 5345 1374
rect -5441 -1278 -5407 1278
rect 5407 -1278 5441 1278
rect -5345 -1374 5345 -1340
<< poly >>
rect -5284 1272 -5218 1288
rect -5284 1238 -5268 1272
rect -5234 1238 -5218 1272
rect -5284 1222 -5218 1238
rect -5166 1272 -5100 1288
rect -5166 1238 -5150 1272
rect -5116 1238 -5100 1272
rect -5166 1222 -5100 1238
rect -5048 1272 -4982 1288
rect -5048 1238 -5032 1272
rect -4998 1238 -4982 1272
rect -5048 1222 -4982 1238
rect -4930 1272 -4864 1288
rect -4930 1238 -4914 1272
rect -4880 1238 -4864 1272
rect -4930 1222 -4864 1238
rect -4812 1272 -4746 1288
rect -4812 1238 -4796 1272
rect -4762 1238 -4746 1272
rect -4812 1222 -4746 1238
rect -4694 1272 -4628 1288
rect -4694 1238 -4678 1272
rect -4644 1238 -4628 1272
rect -4694 1222 -4628 1238
rect -4576 1272 -4510 1288
rect -4576 1238 -4560 1272
rect -4526 1238 -4510 1272
rect -4576 1222 -4510 1238
rect -4458 1272 -4392 1288
rect -4458 1238 -4442 1272
rect -4408 1238 -4392 1272
rect -4458 1222 -4392 1238
rect -4340 1272 -4274 1288
rect -4340 1238 -4324 1272
rect -4290 1238 -4274 1272
rect -4340 1222 -4274 1238
rect -4222 1272 -4156 1288
rect -4222 1238 -4206 1272
rect -4172 1238 -4156 1272
rect -4222 1222 -4156 1238
rect -4104 1272 -4038 1288
rect -4104 1238 -4088 1272
rect -4054 1238 -4038 1272
rect -4104 1222 -4038 1238
rect -3986 1272 -3920 1288
rect -3986 1238 -3970 1272
rect -3936 1238 -3920 1272
rect -3986 1222 -3920 1238
rect -3868 1272 -3802 1288
rect -3868 1238 -3852 1272
rect -3818 1238 -3802 1272
rect -3868 1222 -3802 1238
rect -3750 1272 -3684 1288
rect -3750 1238 -3734 1272
rect -3700 1238 -3684 1272
rect -3750 1222 -3684 1238
rect -3632 1272 -3566 1288
rect -3632 1238 -3616 1272
rect -3582 1238 -3566 1272
rect -3632 1222 -3566 1238
rect -3514 1272 -3448 1288
rect -3514 1238 -3498 1272
rect -3464 1238 -3448 1272
rect -3514 1222 -3448 1238
rect -3396 1272 -3330 1288
rect -3396 1238 -3380 1272
rect -3346 1238 -3330 1272
rect -3396 1222 -3330 1238
rect -3278 1272 -3212 1288
rect -3278 1238 -3262 1272
rect -3228 1238 -3212 1272
rect -3278 1222 -3212 1238
rect -3160 1272 -3094 1288
rect -3160 1238 -3144 1272
rect -3110 1238 -3094 1272
rect -3160 1222 -3094 1238
rect -3042 1272 -2976 1288
rect -3042 1238 -3026 1272
rect -2992 1238 -2976 1272
rect -3042 1222 -2976 1238
rect -2924 1272 -2858 1288
rect -2924 1238 -2908 1272
rect -2874 1238 -2858 1272
rect -2924 1222 -2858 1238
rect -2806 1272 -2740 1288
rect -2806 1238 -2790 1272
rect -2756 1238 -2740 1272
rect -2806 1222 -2740 1238
rect -2688 1272 -2622 1288
rect -2688 1238 -2672 1272
rect -2638 1238 -2622 1272
rect -2688 1222 -2622 1238
rect -2570 1272 -2504 1288
rect -2570 1238 -2554 1272
rect -2520 1238 -2504 1272
rect -2570 1222 -2504 1238
rect -2452 1272 -2386 1288
rect -2452 1238 -2436 1272
rect -2402 1238 -2386 1272
rect -2452 1222 -2386 1238
rect -2334 1272 -2268 1288
rect -2334 1238 -2318 1272
rect -2284 1238 -2268 1272
rect -2334 1222 -2268 1238
rect -2216 1272 -2150 1288
rect -2216 1238 -2200 1272
rect -2166 1238 -2150 1272
rect -2216 1222 -2150 1238
rect -2098 1272 -2032 1288
rect -2098 1238 -2082 1272
rect -2048 1238 -2032 1272
rect -2098 1222 -2032 1238
rect -1980 1272 -1914 1288
rect -1980 1238 -1964 1272
rect -1930 1238 -1914 1272
rect -1980 1222 -1914 1238
rect -1862 1272 -1796 1288
rect -1862 1238 -1846 1272
rect -1812 1238 -1796 1272
rect -1862 1222 -1796 1238
rect -1744 1272 -1678 1288
rect -1744 1238 -1728 1272
rect -1694 1238 -1678 1272
rect -1744 1222 -1678 1238
rect -1626 1272 -1560 1288
rect -1626 1238 -1610 1272
rect -1576 1238 -1560 1272
rect -1626 1222 -1560 1238
rect -1508 1272 -1442 1288
rect -1508 1238 -1492 1272
rect -1458 1238 -1442 1272
rect -1508 1222 -1442 1238
rect -1390 1272 -1324 1288
rect -1390 1238 -1374 1272
rect -1340 1238 -1324 1272
rect -1390 1222 -1324 1238
rect -1272 1272 -1206 1288
rect -1272 1238 -1256 1272
rect -1222 1238 -1206 1272
rect -1272 1222 -1206 1238
rect -1154 1272 -1088 1288
rect -1154 1238 -1138 1272
rect -1104 1238 -1088 1272
rect -1154 1222 -1088 1238
rect -1036 1272 -970 1288
rect -1036 1238 -1020 1272
rect -986 1238 -970 1272
rect -1036 1222 -970 1238
rect -918 1272 -852 1288
rect -918 1238 -902 1272
rect -868 1238 -852 1272
rect -918 1222 -852 1238
rect -800 1272 -734 1288
rect -800 1238 -784 1272
rect -750 1238 -734 1272
rect -800 1222 -734 1238
rect -682 1272 -616 1288
rect -682 1238 -666 1272
rect -632 1238 -616 1272
rect -682 1222 -616 1238
rect -564 1272 -498 1288
rect -564 1238 -548 1272
rect -514 1238 -498 1272
rect -564 1222 -498 1238
rect -446 1272 -380 1288
rect -446 1238 -430 1272
rect -396 1238 -380 1272
rect -446 1222 -380 1238
rect -328 1272 -262 1288
rect -328 1238 -312 1272
rect -278 1238 -262 1272
rect -328 1222 -262 1238
rect -210 1272 -144 1288
rect -210 1238 -194 1272
rect -160 1238 -144 1272
rect -210 1222 -144 1238
rect -92 1272 -26 1288
rect -92 1238 -76 1272
rect -42 1238 -26 1272
rect -92 1222 -26 1238
rect 26 1272 92 1288
rect 26 1238 42 1272
rect 76 1238 92 1272
rect 26 1222 92 1238
rect 144 1272 210 1288
rect 144 1238 160 1272
rect 194 1238 210 1272
rect 144 1222 210 1238
rect 262 1272 328 1288
rect 262 1238 278 1272
rect 312 1238 328 1272
rect 262 1222 328 1238
rect 380 1272 446 1288
rect 380 1238 396 1272
rect 430 1238 446 1272
rect 380 1222 446 1238
rect 498 1272 564 1288
rect 498 1238 514 1272
rect 548 1238 564 1272
rect 498 1222 564 1238
rect 616 1272 682 1288
rect 616 1238 632 1272
rect 666 1238 682 1272
rect 616 1222 682 1238
rect 734 1272 800 1288
rect 734 1238 750 1272
rect 784 1238 800 1272
rect 734 1222 800 1238
rect 852 1272 918 1288
rect 852 1238 868 1272
rect 902 1238 918 1272
rect 852 1222 918 1238
rect 970 1272 1036 1288
rect 970 1238 986 1272
rect 1020 1238 1036 1272
rect 970 1222 1036 1238
rect 1088 1272 1154 1288
rect 1088 1238 1104 1272
rect 1138 1238 1154 1272
rect 1088 1222 1154 1238
rect 1206 1272 1272 1288
rect 1206 1238 1222 1272
rect 1256 1238 1272 1272
rect 1206 1222 1272 1238
rect 1324 1272 1390 1288
rect 1324 1238 1340 1272
rect 1374 1238 1390 1272
rect 1324 1222 1390 1238
rect 1442 1272 1508 1288
rect 1442 1238 1458 1272
rect 1492 1238 1508 1272
rect 1442 1222 1508 1238
rect 1560 1272 1626 1288
rect 1560 1238 1576 1272
rect 1610 1238 1626 1272
rect 1560 1222 1626 1238
rect 1678 1272 1744 1288
rect 1678 1238 1694 1272
rect 1728 1238 1744 1272
rect 1678 1222 1744 1238
rect 1796 1272 1862 1288
rect 1796 1238 1812 1272
rect 1846 1238 1862 1272
rect 1796 1222 1862 1238
rect 1914 1272 1980 1288
rect 1914 1238 1930 1272
rect 1964 1238 1980 1272
rect 1914 1222 1980 1238
rect 2032 1272 2098 1288
rect 2032 1238 2048 1272
rect 2082 1238 2098 1272
rect 2032 1222 2098 1238
rect 2150 1272 2216 1288
rect 2150 1238 2166 1272
rect 2200 1238 2216 1272
rect 2150 1222 2216 1238
rect 2268 1272 2334 1288
rect 2268 1238 2284 1272
rect 2318 1238 2334 1272
rect 2268 1222 2334 1238
rect 2386 1272 2452 1288
rect 2386 1238 2402 1272
rect 2436 1238 2452 1272
rect 2386 1222 2452 1238
rect 2504 1272 2570 1288
rect 2504 1238 2520 1272
rect 2554 1238 2570 1272
rect 2504 1222 2570 1238
rect 2622 1272 2688 1288
rect 2622 1238 2638 1272
rect 2672 1238 2688 1272
rect 2622 1222 2688 1238
rect 2740 1272 2806 1288
rect 2740 1238 2756 1272
rect 2790 1238 2806 1272
rect 2740 1222 2806 1238
rect 2858 1272 2924 1288
rect 2858 1238 2874 1272
rect 2908 1238 2924 1272
rect 2858 1222 2924 1238
rect 2976 1272 3042 1288
rect 2976 1238 2992 1272
rect 3026 1238 3042 1272
rect 2976 1222 3042 1238
rect 3094 1272 3160 1288
rect 3094 1238 3110 1272
rect 3144 1238 3160 1272
rect 3094 1222 3160 1238
rect 3212 1272 3278 1288
rect 3212 1238 3228 1272
rect 3262 1238 3278 1272
rect 3212 1222 3278 1238
rect 3330 1272 3396 1288
rect 3330 1238 3346 1272
rect 3380 1238 3396 1272
rect 3330 1222 3396 1238
rect 3448 1272 3514 1288
rect 3448 1238 3464 1272
rect 3498 1238 3514 1272
rect 3448 1222 3514 1238
rect 3566 1272 3632 1288
rect 3566 1238 3582 1272
rect 3616 1238 3632 1272
rect 3566 1222 3632 1238
rect 3684 1272 3750 1288
rect 3684 1238 3700 1272
rect 3734 1238 3750 1272
rect 3684 1222 3750 1238
rect 3802 1272 3868 1288
rect 3802 1238 3818 1272
rect 3852 1238 3868 1272
rect 3802 1222 3868 1238
rect 3920 1272 3986 1288
rect 3920 1238 3936 1272
rect 3970 1238 3986 1272
rect 3920 1222 3986 1238
rect 4038 1272 4104 1288
rect 4038 1238 4054 1272
rect 4088 1238 4104 1272
rect 4038 1222 4104 1238
rect 4156 1272 4222 1288
rect 4156 1238 4172 1272
rect 4206 1238 4222 1272
rect 4156 1222 4222 1238
rect 4274 1272 4340 1288
rect 4274 1238 4290 1272
rect 4324 1238 4340 1272
rect 4274 1222 4340 1238
rect 4392 1272 4458 1288
rect 4392 1238 4408 1272
rect 4442 1238 4458 1272
rect 4392 1222 4458 1238
rect 4510 1272 4576 1288
rect 4510 1238 4526 1272
rect 4560 1238 4576 1272
rect 4510 1222 4576 1238
rect 4628 1272 4694 1288
rect 4628 1238 4644 1272
rect 4678 1238 4694 1272
rect 4628 1222 4694 1238
rect 4746 1272 4812 1288
rect 4746 1238 4762 1272
rect 4796 1238 4812 1272
rect 4746 1222 4812 1238
rect 4864 1272 4930 1288
rect 4864 1238 4880 1272
rect 4914 1238 4930 1272
rect 4864 1222 4930 1238
rect 4982 1272 5048 1288
rect 4982 1238 4998 1272
rect 5032 1238 5048 1272
rect 4982 1222 5048 1238
rect 5100 1272 5166 1288
rect 5100 1238 5116 1272
rect 5150 1238 5166 1272
rect 5100 1222 5166 1238
rect 5218 1272 5284 1288
rect 5218 1238 5234 1272
rect 5268 1238 5284 1272
rect 5218 1222 5284 1238
rect -5281 1200 -5221 1222
rect -5163 1200 -5103 1222
rect -5045 1200 -4985 1222
rect -4927 1200 -4867 1222
rect -4809 1200 -4749 1222
rect -4691 1200 -4631 1222
rect -4573 1200 -4513 1222
rect -4455 1200 -4395 1222
rect -4337 1200 -4277 1222
rect -4219 1200 -4159 1222
rect -4101 1200 -4041 1222
rect -3983 1200 -3923 1222
rect -3865 1200 -3805 1222
rect -3747 1200 -3687 1222
rect -3629 1200 -3569 1222
rect -3511 1200 -3451 1222
rect -3393 1200 -3333 1222
rect -3275 1200 -3215 1222
rect -3157 1200 -3097 1222
rect -3039 1200 -2979 1222
rect -2921 1200 -2861 1222
rect -2803 1200 -2743 1222
rect -2685 1200 -2625 1222
rect -2567 1200 -2507 1222
rect -2449 1200 -2389 1222
rect -2331 1200 -2271 1222
rect -2213 1200 -2153 1222
rect -2095 1200 -2035 1222
rect -1977 1200 -1917 1222
rect -1859 1200 -1799 1222
rect -1741 1200 -1681 1222
rect -1623 1200 -1563 1222
rect -1505 1200 -1445 1222
rect -1387 1200 -1327 1222
rect -1269 1200 -1209 1222
rect -1151 1200 -1091 1222
rect -1033 1200 -973 1222
rect -915 1200 -855 1222
rect -797 1200 -737 1222
rect -679 1200 -619 1222
rect -561 1200 -501 1222
rect -443 1200 -383 1222
rect -325 1200 -265 1222
rect -207 1200 -147 1222
rect -89 1200 -29 1222
rect 29 1200 89 1222
rect 147 1200 207 1222
rect 265 1200 325 1222
rect 383 1200 443 1222
rect 501 1200 561 1222
rect 619 1200 679 1222
rect 737 1200 797 1222
rect 855 1200 915 1222
rect 973 1200 1033 1222
rect 1091 1200 1151 1222
rect 1209 1200 1269 1222
rect 1327 1200 1387 1222
rect 1445 1200 1505 1222
rect 1563 1200 1623 1222
rect 1681 1200 1741 1222
rect 1799 1200 1859 1222
rect 1917 1200 1977 1222
rect 2035 1200 2095 1222
rect 2153 1200 2213 1222
rect 2271 1200 2331 1222
rect 2389 1200 2449 1222
rect 2507 1200 2567 1222
rect 2625 1200 2685 1222
rect 2743 1200 2803 1222
rect 2861 1200 2921 1222
rect 2979 1200 3039 1222
rect 3097 1200 3157 1222
rect 3215 1200 3275 1222
rect 3333 1200 3393 1222
rect 3451 1200 3511 1222
rect 3569 1200 3629 1222
rect 3687 1200 3747 1222
rect 3805 1200 3865 1222
rect 3923 1200 3983 1222
rect 4041 1200 4101 1222
rect 4159 1200 4219 1222
rect 4277 1200 4337 1222
rect 4395 1200 4455 1222
rect 4513 1200 4573 1222
rect 4631 1200 4691 1222
rect 4749 1200 4809 1222
rect 4867 1200 4927 1222
rect 4985 1200 5045 1222
rect 5103 1200 5163 1222
rect 5221 1200 5281 1222
rect -5281 -1222 -5221 -1200
rect -5163 -1222 -5103 -1200
rect -5045 -1222 -4985 -1200
rect -4927 -1222 -4867 -1200
rect -4809 -1222 -4749 -1200
rect -4691 -1222 -4631 -1200
rect -4573 -1222 -4513 -1200
rect -4455 -1222 -4395 -1200
rect -4337 -1222 -4277 -1200
rect -4219 -1222 -4159 -1200
rect -4101 -1222 -4041 -1200
rect -3983 -1222 -3923 -1200
rect -3865 -1222 -3805 -1200
rect -3747 -1222 -3687 -1200
rect -3629 -1222 -3569 -1200
rect -3511 -1222 -3451 -1200
rect -3393 -1222 -3333 -1200
rect -3275 -1222 -3215 -1200
rect -3157 -1222 -3097 -1200
rect -3039 -1222 -2979 -1200
rect -2921 -1222 -2861 -1200
rect -2803 -1222 -2743 -1200
rect -2685 -1222 -2625 -1200
rect -2567 -1222 -2507 -1200
rect -2449 -1222 -2389 -1200
rect -2331 -1222 -2271 -1200
rect -2213 -1222 -2153 -1200
rect -2095 -1222 -2035 -1200
rect -1977 -1222 -1917 -1200
rect -1859 -1222 -1799 -1200
rect -1741 -1222 -1681 -1200
rect -1623 -1222 -1563 -1200
rect -1505 -1222 -1445 -1200
rect -1387 -1222 -1327 -1200
rect -1269 -1222 -1209 -1200
rect -1151 -1222 -1091 -1200
rect -1033 -1222 -973 -1200
rect -915 -1222 -855 -1200
rect -797 -1222 -737 -1200
rect -679 -1222 -619 -1200
rect -561 -1222 -501 -1200
rect -443 -1222 -383 -1200
rect -325 -1222 -265 -1200
rect -207 -1222 -147 -1200
rect -89 -1222 -29 -1200
rect 29 -1222 89 -1200
rect 147 -1222 207 -1200
rect 265 -1222 325 -1200
rect 383 -1222 443 -1200
rect 501 -1222 561 -1200
rect 619 -1222 679 -1200
rect 737 -1222 797 -1200
rect 855 -1222 915 -1200
rect 973 -1222 1033 -1200
rect 1091 -1222 1151 -1200
rect 1209 -1222 1269 -1200
rect 1327 -1222 1387 -1200
rect 1445 -1222 1505 -1200
rect 1563 -1222 1623 -1200
rect 1681 -1222 1741 -1200
rect 1799 -1222 1859 -1200
rect 1917 -1222 1977 -1200
rect 2035 -1222 2095 -1200
rect 2153 -1222 2213 -1200
rect 2271 -1222 2331 -1200
rect 2389 -1222 2449 -1200
rect 2507 -1222 2567 -1200
rect 2625 -1222 2685 -1200
rect 2743 -1222 2803 -1200
rect 2861 -1222 2921 -1200
rect 2979 -1222 3039 -1200
rect 3097 -1222 3157 -1200
rect 3215 -1222 3275 -1200
rect 3333 -1222 3393 -1200
rect 3451 -1222 3511 -1200
rect 3569 -1222 3629 -1200
rect 3687 -1222 3747 -1200
rect 3805 -1222 3865 -1200
rect 3923 -1222 3983 -1200
rect 4041 -1222 4101 -1200
rect 4159 -1222 4219 -1200
rect 4277 -1222 4337 -1200
rect 4395 -1222 4455 -1200
rect 4513 -1222 4573 -1200
rect 4631 -1222 4691 -1200
rect 4749 -1222 4809 -1200
rect 4867 -1222 4927 -1200
rect 4985 -1222 5045 -1200
rect 5103 -1222 5163 -1200
rect 5221 -1222 5281 -1200
rect -5284 -1238 -5218 -1222
rect -5284 -1272 -5268 -1238
rect -5234 -1272 -5218 -1238
rect -5284 -1288 -5218 -1272
rect -5166 -1238 -5100 -1222
rect -5166 -1272 -5150 -1238
rect -5116 -1272 -5100 -1238
rect -5166 -1288 -5100 -1272
rect -5048 -1238 -4982 -1222
rect -5048 -1272 -5032 -1238
rect -4998 -1272 -4982 -1238
rect -5048 -1288 -4982 -1272
rect -4930 -1238 -4864 -1222
rect -4930 -1272 -4914 -1238
rect -4880 -1272 -4864 -1238
rect -4930 -1288 -4864 -1272
rect -4812 -1238 -4746 -1222
rect -4812 -1272 -4796 -1238
rect -4762 -1272 -4746 -1238
rect -4812 -1288 -4746 -1272
rect -4694 -1238 -4628 -1222
rect -4694 -1272 -4678 -1238
rect -4644 -1272 -4628 -1238
rect -4694 -1288 -4628 -1272
rect -4576 -1238 -4510 -1222
rect -4576 -1272 -4560 -1238
rect -4526 -1272 -4510 -1238
rect -4576 -1288 -4510 -1272
rect -4458 -1238 -4392 -1222
rect -4458 -1272 -4442 -1238
rect -4408 -1272 -4392 -1238
rect -4458 -1288 -4392 -1272
rect -4340 -1238 -4274 -1222
rect -4340 -1272 -4324 -1238
rect -4290 -1272 -4274 -1238
rect -4340 -1288 -4274 -1272
rect -4222 -1238 -4156 -1222
rect -4222 -1272 -4206 -1238
rect -4172 -1272 -4156 -1238
rect -4222 -1288 -4156 -1272
rect -4104 -1238 -4038 -1222
rect -4104 -1272 -4088 -1238
rect -4054 -1272 -4038 -1238
rect -4104 -1288 -4038 -1272
rect -3986 -1238 -3920 -1222
rect -3986 -1272 -3970 -1238
rect -3936 -1272 -3920 -1238
rect -3986 -1288 -3920 -1272
rect -3868 -1238 -3802 -1222
rect -3868 -1272 -3852 -1238
rect -3818 -1272 -3802 -1238
rect -3868 -1288 -3802 -1272
rect -3750 -1238 -3684 -1222
rect -3750 -1272 -3734 -1238
rect -3700 -1272 -3684 -1238
rect -3750 -1288 -3684 -1272
rect -3632 -1238 -3566 -1222
rect -3632 -1272 -3616 -1238
rect -3582 -1272 -3566 -1238
rect -3632 -1288 -3566 -1272
rect -3514 -1238 -3448 -1222
rect -3514 -1272 -3498 -1238
rect -3464 -1272 -3448 -1238
rect -3514 -1288 -3448 -1272
rect -3396 -1238 -3330 -1222
rect -3396 -1272 -3380 -1238
rect -3346 -1272 -3330 -1238
rect -3396 -1288 -3330 -1272
rect -3278 -1238 -3212 -1222
rect -3278 -1272 -3262 -1238
rect -3228 -1272 -3212 -1238
rect -3278 -1288 -3212 -1272
rect -3160 -1238 -3094 -1222
rect -3160 -1272 -3144 -1238
rect -3110 -1272 -3094 -1238
rect -3160 -1288 -3094 -1272
rect -3042 -1238 -2976 -1222
rect -3042 -1272 -3026 -1238
rect -2992 -1272 -2976 -1238
rect -3042 -1288 -2976 -1272
rect -2924 -1238 -2858 -1222
rect -2924 -1272 -2908 -1238
rect -2874 -1272 -2858 -1238
rect -2924 -1288 -2858 -1272
rect -2806 -1238 -2740 -1222
rect -2806 -1272 -2790 -1238
rect -2756 -1272 -2740 -1238
rect -2806 -1288 -2740 -1272
rect -2688 -1238 -2622 -1222
rect -2688 -1272 -2672 -1238
rect -2638 -1272 -2622 -1238
rect -2688 -1288 -2622 -1272
rect -2570 -1238 -2504 -1222
rect -2570 -1272 -2554 -1238
rect -2520 -1272 -2504 -1238
rect -2570 -1288 -2504 -1272
rect -2452 -1238 -2386 -1222
rect -2452 -1272 -2436 -1238
rect -2402 -1272 -2386 -1238
rect -2452 -1288 -2386 -1272
rect -2334 -1238 -2268 -1222
rect -2334 -1272 -2318 -1238
rect -2284 -1272 -2268 -1238
rect -2334 -1288 -2268 -1272
rect -2216 -1238 -2150 -1222
rect -2216 -1272 -2200 -1238
rect -2166 -1272 -2150 -1238
rect -2216 -1288 -2150 -1272
rect -2098 -1238 -2032 -1222
rect -2098 -1272 -2082 -1238
rect -2048 -1272 -2032 -1238
rect -2098 -1288 -2032 -1272
rect -1980 -1238 -1914 -1222
rect -1980 -1272 -1964 -1238
rect -1930 -1272 -1914 -1238
rect -1980 -1288 -1914 -1272
rect -1862 -1238 -1796 -1222
rect -1862 -1272 -1846 -1238
rect -1812 -1272 -1796 -1238
rect -1862 -1288 -1796 -1272
rect -1744 -1238 -1678 -1222
rect -1744 -1272 -1728 -1238
rect -1694 -1272 -1678 -1238
rect -1744 -1288 -1678 -1272
rect -1626 -1238 -1560 -1222
rect -1626 -1272 -1610 -1238
rect -1576 -1272 -1560 -1238
rect -1626 -1288 -1560 -1272
rect -1508 -1238 -1442 -1222
rect -1508 -1272 -1492 -1238
rect -1458 -1272 -1442 -1238
rect -1508 -1288 -1442 -1272
rect -1390 -1238 -1324 -1222
rect -1390 -1272 -1374 -1238
rect -1340 -1272 -1324 -1238
rect -1390 -1288 -1324 -1272
rect -1272 -1238 -1206 -1222
rect -1272 -1272 -1256 -1238
rect -1222 -1272 -1206 -1238
rect -1272 -1288 -1206 -1272
rect -1154 -1238 -1088 -1222
rect -1154 -1272 -1138 -1238
rect -1104 -1272 -1088 -1238
rect -1154 -1288 -1088 -1272
rect -1036 -1238 -970 -1222
rect -1036 -1272 -1020 -1238
rect -986 -1272 -970 -1238
rect -1036 -1288 -970 -1272
rect -918 -1238 -852 -1222
rect -918 -1272 -902 -1238
rect -868 -1272 -852 -1238
rect -918 -1288 -852 -1272
rect -800 -1238 -734 -1222
rect -800 -1272 -784 -1238
rect -750 -1272 -734 -1238
rect -800 -1288 -734 -1272
rect -682 -1238 -616 -1222
rect -682 -1272 -666 -1238
rect -632 -1272 -616 -1238
rect -682 -1288 -616 -1272
rect -564 -1238 -498 -1222
rect -564 -1272 -548 -1238
rect -514 -1272 -498 -1238
rect -564 -1288 -498 -1272
rect -446 -1238 -380 -1222
rect -446 -1272 -430 -1238
rect -396 -1272 -380 -1238
rect -446 -1288 -380 -1272
rect -328 -1238 -262 -1222
rect -328 -1272 -312 -1238
rect -278 -1272 -262 -1238
rect -328 -1288 -262 -1272
rect -210 -1238 -144 -1222
rect -210 -1272 -194 -1238
rect -160 -1272 -144 -1238
rect -210 -1288 -144 -1272
rect -92 -1238 -26 -1222
rect -92 -1272 -76 -1238
rect -42 -1272 -26 -1238
rect -92 -1288 -26 -1272
rect 26 -1238 92 -1222
rect 26 -1272 42 -1238
rect 76 -1272 92 -1238
rect 26 -1288 92 -1272
rect 144 -1238 210 -1222
rect 144 -1272 160 -1238
rect 194 -1272 210 -1238
rect 144 -1288 210 -1272
rect 262 -1238 328 -1222
rect 262 -1272 278 -1238
rect 312 -1272 328 -1238
rect 262 -1288 328 -1272
rect 380 -1238 446 -1222
rect 380 -1272 396 -1238
rect 430 -1272 446 -1238
rect 380 -1288 446 -1272
rect 498 -1238 564 -1222
rect 498 -1272 514 -1238
rect 548 -1272 564 -1238
rect 498 -1288 564 -1272
rect 616 -1238 682 -1222
rect 616 -1272 632 -1238
rect 666 -1272 682 -1238
rect 616 -1288 682 -1272
rect 734 -1238 800 -1222
rect 734 -1272 750 -1238
rect 784 -1272 800 -1238
rect 734 -1288 800 -1272
rect 852 -1238 918 -1222
rect 852 -1272 868 -1238
rect 902 -1272 918 -1238
rect 852 -1288 918 -1272
rect 970 -1238 1036 -1222
rect 970 -1272 986 -1238
rect 1020 -1272 1036 -1238
rect 970 -1288 1036 -1272
rect 1088 -1238 1154 -1222
rect 1088 -1272 1104 -1238
rect 1138 -1272 1154 -1238
rect 1088 -1288 1154 -1272
rect 1206 -1238 1272 -1222
rect 1206 -1272 1222 -1238
rect 1256 -1272 1272 -1238
rect 1206 -1288 1272 -1272
rect 1324 -1238 1390 -1222
rect 1324 -1272 1340 -1238
rect 1374 -1272 1390 -1238
rect 1324 -1288 1390 -1272
rect 1442 -1238 1508 -1222
rect 1442 -1272 1458 -1238
rect 1492 -1272 1508 -1238
rect 1442 -1288 1508 -1272
rect 1560 -1238 1626 -1222
rect 1560 -1272 1576 -1238
rect 1610 -1272 1626 -1238
rect 1560 -1288 1626 -1272
rect 1678 -1238 1744 -1222
rect 1678 -1272 1694 -1238
rect 1728 -1272 1744 -1238
rect 1678 -1288 1744 -1272
rect 1796 -1238 1862 -1222
rect 1796 -1272 1812 -1238
rect 1846 -1272 1862 -1238
rect 1796 -1288 1862 -1272
rect 1914 -1238 1980 -1222
rect 1914 -1272 1930 -1238
rect 1964 -1272 1980 -1238
rect 1914 -1288 1980 -1272
rect 2032 -1238 2098 -1222
rect 2032 -1272 2048 -1238
rect 2082 -1272 2098 -1238
rect 2032 -1288 2098 -1272
rect 2150 -1238 2216 -1222
rect 2150 -1272 2166 -1238
rect 2200 -1272 2216 -1238
rect 2150 -1288 2216 -1272
rect 2268 -1238 2334 -1222
rect 2268 -1272 2284 -1238
rect 2318 -1272 2334 -1238
rect 2268 -1288 2334 -1272
rect 2386 -1238 2452 -1222
rect 2386 -1272 2402 -1238
rect 2436 -1272 2452 -1238
rect 2386 -1288 2452 -1272
rect 2504 -1238 2570 -1222
rect 2504 -1272 2520 -1238
rect 2554 -1272 2570 -1238
rect 2504 -1288 2570 -1272
rect 2622 -1238 2688 -1222
rect 2622 -1272 2638 -1238
rect 2672 -1272 2688 -1238
rect 2622 -1288 2688 -1272
rect 2740 -1238 2806 -1222
rect 2740 -1272 2756 -1238
rect 2790 -1272 2806 -1238
rect 2740 -1288 2806 -1272
rect 2858 -1238 2924 -1222
rect 2858 -1272 2874 -1238
rect 2908 -1272 2924 -1238
rect 2858 -1288 2924 -1272
rect 2976 -1238 3042 -1222
rect 2976 -1272 2992 -1238
rect 3026 -1272 3042 -1238
rect 2976 -1288 3042 -1272
rect 3094 -1238 3160 -1222
rect 3094 -1272 3110 -1238
rect 3144 -1272 3160 -1238
rect 3094 -1288 3160 -1272
rect 3212 -1238 3278 -1222
rect 3212 -1272 3228 -1238
rect 3262 -1272 3278 -1238
rect 3212 -1288 3278 -1272
rect 3330 -1238 3396 -1222
rect 3330 -1272 3346 -1238
rect 3380 -1272 3396 -1238
rect 3330 -1288 3396 -1272
rect 3448 -1238 3514 -1222
rect 3448 -1272 3464 -1238
rect 3498 -1272 3514 -1238
rect 3448 -1288 3514 -1272
rect 3566 -1238 3632 -1222
rect 3566 -1272 3582 -1238
rect 3616 -1272 3632 -1238
rect 3566 -1288 3632 -1272
rect 3684 -1238 3750 -1222
rect 3684 -1272 3700 -1238
rect 3734 -1272 3750 -1238
rect 3684 -1288 3750 -1272
rect 3802 -1238 3868 -1222
rect 3802 -1272 3818 -1238
rect 3852 -1272 3868 -1238
rect 3802 -1288 3868 -1272
rect 3920 -1238 3986 -1222
rect 3920 -1272 3936 -1238
rect 3970 -1272 3986 -1238
rect 3920 -1288 3986 -1272
rect 4038 -1238 4104 -1222
rect 4038 -1272 4054 -1238
rect 4088 -1272 4104 -1238
rect 4038 -1288 4104 -1272
rect 4156 -1238 4222 -1222
rect 4156 -1272 4172 -1238
rect 4206 -1272 4222 -1238
rect 4156 -1288 4222 -1272
rect 4274 -1238 4340 -1222
rect 4274 -1272 4290 -1238
rect 4324 -1272 4340 -1238
rect 4274 -1288 4340 -1272
rect 4392 -1238 4458 -1222
rect 4392 -1272 4408 -1238
rect 4442 -1272 4458 -1238
rect 4392 -1288 4458 -1272
rect 4510 -1238 4576 -1222
rect 4510 -1272 4526 -1238
rect 4560 -1272 4576 -1238
rect 4510 -1288 4576 -1272
rect 4628 -1238 4694 -1222
rect 4628 -1272 4644 -1238
rect 4678 -1272 4694 -1238
rect 4628 -1288 4694 -1272
rect 4746 -1238 4812 -1222
rect 4746 -1272 4762 -1238
rect 4796 -1272 4812 -1238
rect 4746 -1288 4812 -1272
rect 4864 -1238 4930 -1222
rect 4864 -1272 4880 -1238
rect 4914 -1272 4930 -1238
rect 4864 -1288 4930 -1272
rect 4982 -1238 5048 -1222
rect 4982 -1272 4998 -1238
rect 5032 -1272 5048 -1238
rect 4982 -1288 5048 -1272
rect 5100 -1238 5166 -1222
rect 5100 -1272 5116 -1238
rect 5150 -1272 5166 -1238
rect 5100 -1288 5166 -1272
rect 5218 -1238 5284 -1222
rect 5218 -1272 5234 -1238
rect 5268 -1272 5284 -1238
rect 5218 -1288 5284 -1272
<< polycont >>
rect -5268 1238 -5234 1272
rect -5150 1238 -5116 1272
rect -5032 1238 -4998 1272
rect -4914 1238 -4880 1272
rect -4796 1238 -4762 1272
rect -4678 1238 -4644 1272
rect -4560 1238 -4526 1272
rect -4442 1238 -4408 1272
rect -4324 1238 -4290 1272
rect -4206 1238 -4172 1272
rect -4088 1238 -4054 1272
rect -3970 1238 -3936 1272
rect -3852 1238 -3818 1272
rect -3734 1238 -3700 1272
rect -3616 1238 -3582 1272
rect -3498 1238 -3464 1272
rect -3380 1238 -3346 1272
rect -3262 1238 -3228 1272
rect -3144 1238 -3110 1272
rect -3026 1238 -2992 1272
rect -2908 1238 -2874 1272
rect -2790 1238 -2756 1272
rect -2672 1238 -2638 1272
rect -2554 1238 -2520 1272
rect -2436 1238 -2402 1272
rect -2318 1238 -2284 1272
rect -2200 1238 -2166 1272
rect -2082 1238 -2048 1272
rect -1964 1238 -1930 1272
rect -1846 1238 -1812 1272
rect -1728 1238 -1694 1272
rect -1610 1238 -1576 1272
rect -1492 1238 -1458 1272
rect -1374 1238 -1340 1272
rect -1256 1238 -1222 1272
rect -1138 1238 -1104 1272
rect -1020 1238 -986 1272
rect -902 1238 -868 1272
rect -784 1238 -750 1272
rect -666 1238 -632 1272
rect -548 1238 -514 1272
rect -430 1238 -396 1272
rect -312 1238 -278 1272
rect -194 1238 -160 1272
rect -76 1238 -42 1272
rect 42 1238 76 1272
rect 160 1238 194 1272
rect 278 1238 312 1272
rect 396 1238 430 1272
rect 514 1238 548 1272
rect 632 1238 666 1272
rect 750 1238 784 1272
rect 868 1238 902 1272
rect 986 1238 1020 1272
rect 1104 1238 1138 1272
rect 1222 1238 1256 1272
rect 1340 1238 1374 1272
rect 1458 1238 1492 1272
rect 1576 1238 1610 1272
rect 1694 1238 1728 1272
rect 1812 1238 1846 1272
rect 1930 1238 1964 1272
rect 2048 1238 2082 1272
rect 2166 1238 2200 1272
rect 2284 1238 2318 1272
rect 2402 1238 2436 1272
rect 2520 1238 2554 1272
rect 2638 1238 2672 1272
rect 2756 1238 2790 1272
rect 2874 1238 2908 1272
rect 2992 1238 3026 1272
rect 3110 1238 3144 1272
rect 3228 1238 3262 1272
rect 3346 1238 3380 1272
rect 3464 1238 3498 1272
rect 3582 1238 3616 1272
rect 3700 1238 3734 1272
rect 3818 1238 3852 1272
rect 3936 1238 3970 1272
rect 4054 1238 4088 1272
rect 4172 1238 4206 1272
rect 4290 1238 4324 1272
rect 4408 1238 4442 1272
rect 4526 1238 4560 1272
rect 4644 1238 4678 1272
rect 4762 1238 4796 1272
rect 4880 1238 4914 1272
rect 4998 1238 5032 1272
rect 5116 1238 5150 1272
rect 5234 1238 5268 1272
rect -5268 -1272 -5234 -1238
rect -5150 -1272 -5116 -1238
rect -5032 -1272 -4998 -1238
rect -4914 -1272 -4880 -1238
rect -4796 -1272 -4762 -1238
rect -4678 -1272 -4644 -1238
rect -4560 -1272 -4526 -1238
rect -4442 -1272 -4408 -1238
rect -4324 -1272 -4290 -1238
rect -4206 -1272 -4172 -1238
rect -4088 -1272 -4054 -1238
rect -3970 -1272 -3936 -1238
rect -3852 -1272 -3818 -1238
rect -3734 -1272 -3700 -1238
rect -3616 -1272 -3582 -1238
rect -3498 -1272 -3464 -1238
rect -3380 -1272 -3346 -1238
rect -3262 -1272 -3228 -1238
rect -3144 -1272 -3110 -1238
rect -3026 -1272 -2992 -1238
rect -2908 -1272 -2874 -1238
rect -2790 -1272 -2756 -1238
rect -2672 -1272 -2638 -1238
rect -2554 -1272 -2520 -1238
rect -2436 -1272 -2402 -1238
rect -2318 -1272 -2284 -1238
rect -2200 -1272 -2166 -1238
rect -2082 -1272 -2048 -1238
rect -1964 -1272 -1930 -1238
rect -1846 -1272 -1812 -1238
rect -1728 -1272 -1694 -1238
rect -1610 -1272 -1576 -1238
rect -1492 -1272 -1458 -1238
rect -1374 -1272 -1340 -1238
rect -1256 -1272 -1222 -1238
rect -1138 -1272 -1104 -1238
rect -1020 -1272 -986 -1238
rect -902 -1272 -868 -1238
rect -784 -1272 -750 -1238
rect -666 -1272 -632 -1238
rect -548 -1272 -514 -1238
rect -430 -1272 -396 -1238
rect -312 -1272 -278 -1238
rect -194 -1272 -160 -1238
rect -76 -1272 -42 -1238
rect 42 -1272 76 -1238
rect 160 -1272 194 -1238
rect 278 -1272 312 -1238
rect 396 -1272 430 -1238
rect 514 -1272 548 -1238
rect 632 -1272 666 -1238
rect 750 -1272 784 -1238
rect 868 -1272 902 -1238
rect 986 -1272 1020 -1238
rect 1104 -1272 1138 -1238
rect 1222 -1272 1256 -1238
rect 1340 -1272 1374 -1238
rect 1458 -1272 1492 -1238
rect 1576 -1272 1610 -1238
rect 1694 -1272 1728 -1238
rect 1812 -1272 1846 -1238
rect 1930 -1272 1964 -1238
rect 2048 -1272 2082 -1238
rect 2166 -1272 2200 -1238
rect 2284 -1272 2318 -1238
rect 2402 -1272 2436 -1238
rect 2520 -1272 2554 -1238
rect 2638 -1272 2672 -1238
rect 2756 -1272 2790 -1238
rect 2874 -1272 2908 -1238
rect 2992 -1272 3026 -1238
rect 3110 -1272 3144 -1238
rect 3228 -1272 3262 -1238
rect 3346 -1272 3380 -1238
rect 3464 -1272 3498 -1238
rect 3582 -1272 3616 -1238
rect 3700 -1272 3734 -1238
rect 3818 -1272 3852 -1238
rect 3936 -1272 3970 -1238
rect 4054 -1272 4088 -1238
rect 4172 -1272 4206 -1238
rect 4290 -1272 4324 -1238
rect 4408 -1272 4442 -1238
rect 4526 -1272 4560 -1238
rect 4644 -1272 4678 -1238
rect 4762 -1272 4796 -1238
rect 4880 -1272 4914 -1238
rect 4998 -1272 5032 -1238
rect 5116 -1272 5150 -1238
rect 5234 -1272 5268 -1238
<< locali >>
rect -5441 1340 -5345 1374
rect 5345 1340 5441 1374
rect -5441 1278 -5407 1340
rect 5407 1278 5441 1340
rect -5284 1238 -5268 1272
rect -5234 1238 -5218 1272
rect -5166 1238 -5150 1272
rect -5116 1238 -5100 1272
rect -5048 1238 -5032 1272
rect -4998 1238 -4982 1272
rect -4930 1238 -4914 1272
rect -4880 1238 -4864 1272
rect -4812 1238 -4796 1272
rect -4762 1238 -4746 1272
rect -4694 1238 -4678 1272
rect -4644 1238 -4628 1272
rect -4576 1238 -4560 1272
rect -4526 1238 -4510 1272
rect -4458 1238 -4442 1272
rect -4408 1238 -4392 1272
rect -4340 1238 -4324 1272
rect -4290 1238 -4274 1272
rect -4222 1238 -4206 1272
rect -4172 1238 -4156 1272
rect -4104 1238 -4088 1272
rect -4054 1238 -4038 1272
rect -3986 1238 -3970 1272
rect -3936 1238 -3920 1272
rect -3868 1238 -3852 1272
rect -3818 1238 -3802 1272
rect -3750 1238 -3734 1272
rect -3700 1238 -3684 1272
rect -3632 1238 -3616 1272
rect -3582 1238 -3566 1272
rect -3514 1238 -3498 1272
rect -3464 1238 -3448 1272
rect -3396 1238 -3380 1272
rect -3346 1238 -3330 1272
rect -3278 1238 -3262 1272
rect -3228 1238 -3212 1272
rect -3160 1238 -3144 1272
rect -3110 1238 -3094 1272
rect -3042 1238 -3026 1272
rect -2992 1238 -2976 1272
rect -2924 1238 -2908 1272
rect -2874 1238 -2858 1272
rect -2806 1238 -2790 1272
rect -2756 1238 -2740 1272
rect -2688 1238 -2672 1272
rect -2638 1238 -2622 1272
rect -2570 1238 -2554 1272
rect -2520 1238 -2504 1272
rect -2452 1238 -2436 1272
rect -2402 1238 -2386 1272
rect -2334 1238 -2318 1272
rect -2284 1238 -2268 1272
rect -2216 1238 -2200 1272
rect -2166 1238 -2150 1272
rect -2098 1238 -2082 1272
rect -2048 1238 -2032 1272
rect -1980 1238 -1964 1272
rect -1930 1238 -1914 1272
rect -1862 1238 -1846 1272
rect -1812 1238 -1796 1272
rect -1744 1238 -1728 1272
rect -1694 1238 -1678 1272
rect -1626 1238 -1610 1272
rect -1576 1238 -1560 1272
rect -1508 1238 -1492 1272
rect -1458 1238 -1442 1272
rect -1390 1238 -1374 1272
rect -1340 1238 -1324 1272
rect -1272 1238 -1256 1272
rect -1222 1238 -1206 1272
rect -1154 1238 -1138 1272
rect -1104 1238 -1088 1272
rect -1036 1238 -1020 1272
rect -986 1238 -970 1272
rect -918 1238 -902 1272
rect -868 1238 -852 1272
rect -800 1238 -784 1272
rect -750 1238 -734 1272
rect -682 1238 -666 1272
rect -632 1238 -616 1272
rect -564 1238 -548 1272
rect -514 1238 -498 1272
rect -446 1238 -430 1272
rect -396 1238 -380 1272
rect -328 1238 -312 1272
rect -278 1238 -262 1272
rect -210 1238 -194 1272
rect -160 1238 -144 1272
rect -92 1238 -76 1272
rect -42 1238 -26 1272
rect 26 1238 42 1272
rect 76 1238 92 1272
rect 144 1238 160 1272
rect 194 1238 210 1272
rect 262 1238 278 1272
rect 312 1238 328 1272
rect 380 1238 396 1272
rect 430 1238 446 1272
rect 498 1238 514 1272
rect 548 1238 564 1272
rect 616 1238 632 1272
rect 666 1238 682 1272
rect 734 1238 750 1272
rect 784 1238 800 1272
rect 852 1238 868 1272
rect 902 1238 918 1272
rect 970 1238 986 1272
rect 1020 1238 1036 1272
rect 1088 1238 1104 1272
rect 1138 1238 1154 1272
rect 1206 1238 1222 1272
rect 1256 1238 1272 1272
rect 1324 1238 1340 1272
rect 1374 1238 1390 1272
rect 1442 1238 1458 1272
rect 1492 1238 1508 1272
rect 1560 1238 1576 1272
rect 1610 1238 1626 1272
rect 1678 1238 1694 1272
rect 1728 1238 1744 1272
rect 1796 1238 1812 1272
rect 1846 1238 1862 1272
rect 1914 1238 1930 1272
rect 1964 1238 1980 1272
rect 2032 1238 2048 1272
rect 2082 1238 2098 1272
rect 2150 1238 2166 1272
rect 2200 1238 2216 1272
rect 2268 1238 2284 1272
rect 2318 1238 2334 1272
rect 2386 1238 2402 1272
rect 2436 1238 2452 1272
rect 2504 1238 2520 1272
rect 2554 1238 2570 1272
rect 2622 1238 2638 1272
rect 2672 1238 2688 1272
rect 2740 1238 2756 1272
rect 2790 1238 2806 1272
rect 2858 1238 2874 1272
rect 2908 1238 2924 1272
rect 2976 1238 2992 1272
rect 3026 1238 3042 1272
rect 3094 1238 3110 1272
rect 3144 1238 3160 1272
rect 3212 1238 3228 1272
rect 3262 1238 3278 1272
rect 3330 1238 3346 1272
rect 3380 1238 3396 1272
rect 3448 1238 3464 1272
rect 3498 1238 3514 1272
rect 3566 1238 3582 1272
rect 3616 1238 3632 1272
rect 3684 1238 3700 1272
rect 3734 1238 3750 1272
rect 3802 1238 3818 1272
rect 3852 1238 3868 1272
rect 3920 1238 3936 1272
rect 3970 1238 3986 1272
rect 4038 1238 4054 1272
rect 4088 1238 4104 1272
rect 4156 1238 4172 1272
rect 4206 1238 4222 1272
rect 4274 1238 4290 1272
rect 4324 1238 4340 1272
rect 4392 1238 4408 1272
rect 4442 1238 4458 1272
rect 4510 1238 4526 1272
rect 4560 1238 4576 1272
rect 4628 1238 4644 1272
rect 4678 1238 4694 1272
rect 4746 1238 4762 1272
rect 4796 1238 4812 1272
rect 4864 1238 4880 1272
rect 4914 1238 4930 1272
rect 4982 1238 4998 1272
rect 5032 1238 5048 1272
rect 5100 1238 5116 1272
rect 5150 1238 5166 1272
rect 5218 1238 5234 1272
rect 5268 1238 5284 1272
rect -5327 1188 -5293 1204
rect -5327 -1204 -5293 -1188
rect -5209 1188 -5175 1204
rect -5209 -1204 -5175 -1188
rect -5091 1188 -5057 1204
rect -5091 -1204 -5057 -1188
rect -4973 1188 -4939 1204
rect -4973 -1204 -4939 -1188
rect -4855 1188 -4821 1204
rect -4855 -1204 -4821 -1188
rect -4737 1188 -4703 1204
rect -4737 -1204 -4703 -1188
rect -4619 1188 -4585 1204
rect -4619 -1204 -4585 -1188
rect -4501 1188 -4467 1204
rect -4501 -1204 -4467 -1188
rect -4383 1188 -4349 1204
rect -4383 -1204 -4349 -1188
rect -4265 1188 -4231 1204
rect -4265 -1204 -4231 -1188
rect -4147 1188 -4113 1204
rect -4147 -1204 -4113 -1188
rect -4029 1188 -3995 1204
rect -4029 -1204 -3995 -1188
rect -3911 1188 -3877 1204
rect -3911 -1204 -3877 -1188
rect -3793 1188 -3759 1204
rect -3793 -1204 -3759 -1188
rect -3675 1188 -3641 1204
rect -3675 -1204 -3641 -1188
rect -3557 1188 -3523 1204
rect -3557 -1204 -3523 -1188
rect -3439 1188 -3405 1204
rect -3439 -1204 -3405 -1188
rect -3321 1188 -3287 1204
rect -3321 -1204 -3287 -1188
rect -3203 1188 -3169 1204
rect -3203 -1204 -3169 -1188
rect -3085 1188 -3051 1204
rect -3085 -1204 -3051 -1188
rect -2967 1188 -2933 1204
rect -2967 -1204 -2933 -1188
rect -2849 1188 -2815 1204
rect -2849 -1204 -2815 -1188
rect -2731 1188 -2697 1204
rect -2731 -1204 -2697 -1188
rect -2613 1188 -2579 1204
rect -2613 -1204 -2579 -1188
rect -2495 1188 -2461 1204
rect -2495 -1204 -2461 -1188
rect -2377 1188 -2343 1204
rect -2377 -1204 -2343 -1188
rect -2259 1188 -2225 1204
rect -2259 -1204 -2225 -1188
rect -2141 1188 -2107 1204
rect -2141 -1204 -2107 -1188
rect -2023 1188 -1989 1204
rect -2023 -1204 -1989 -1188
rect -1905 1188 -1871 1204
rect -1905 -1204 -1871 -1188
rect -1787 1188 -1753 1204
rect -1787 -1204 -1753 -1188
rect -1669 1188 -1635 1204
rect -1669 -1204 -1635 -1188
rect -1551 1188 -1517 1204
rect -1551 -1204 -1517 -1188
rect -1433 1188 -1399 1204
rect -1433 -1204 -1399 -1188
rect -1315 1188 -1281 1204
rect -1315 -1204 -1281 -1188
rect -1197 1188 -1163 1204
rect -1197 -1204 -1163 -1188
rect -1079 1188 -1045 1204
rect -1079 -1204 -1045 -1188
rect -961 1188 -927 1204
rect -961 -1204 -927 -1188
rect -843 1188 -809 1204
rect -843 -1204 -809 -1188
rect -725 1188 -691 1204
rect -725 -1204 -691 -1188
rect -607 1188 -573 1204
rect -607 -1204 -573 -1188
rect -489 1188 -455 1204
rect -489 -1204 -455 -1188
rect -371 1188 -337 1204
rect -371 -1204 -337 -1188
rect -253 1188 -219 1204
rect -253 -1204 -219 -1188
rect -135 1188 -101 1204
rect -135 -1204 -101 -1188
rect -17 1188 17 1204
rect -17 -1204 17 -1188
rect 101 1188 135 1204
rect 101 -1204 135 -1188
rect 219 1188 253 1204
rect 219 -1204 253 -1188
rect 337 1188 371 1204
rect 337 -1204 371 -1188
rect 455 1188 489 1204
rect 455 -1204 489 -1188
rect 573 1188 607 1204
rect 573 -1204 607 -1188
rect 691 1188 725 1204
rect 691 -1204 725 -1188
rect 809 1188 843 1204
rect 809 -1204 843 -1188
rect 927 1188 961 1204
rect 927 -1204 961 -1188
rect 1045 1188 1079 1204
rect 1045 -1204 1079 -1188
rect 1163 1188 1197 1204
rect 1163 -1204 1197 -1188
rect 1281 1188 1315 1204
rect 1281 -1204 1315 -1188
rect 1399 1188 1433 1204
rect 1399 -1204 1433 -1188
rect 1517 1188 1551 1204
rect 1517 -1204 1551 -1188
rect 1635 1188 1669 1204
rect 1635 -1204 1669 -1188
rect 1753 1188 1787 1204
rect 1753 -1204 1787 -1188
rect 1871 1188 1905 1204
rect 1871 -1204 1905 -1188
rect 1989 1188 2023 1204
rect 1989 -1204 2023 -1188
rect 2107 1188 2141 1204
rect 2107 -1204 2141 -1188
rect 2225 1188 2259 1204
rect 2225 -1204 2259 -1188
rect 2343 1188 2377 1204
rect 2343 -1204 2377 -1188
rect 2461 1188 2495 1204
rect 2461 -1204 2495 -1188
rect 2579 1188 2613 1204
rect 2579 -1204 2613 -1188
rect 2697 1188 2731 1204
rect 2697 -1204 2731 -1188
rect 2815 1188 2849 1204
rect 2815 -1204 2849 -1188
rect 2933 1188 2967 1204
rect 2933 -1204 2967 -1188
rect 3051 1188 3085 1204
rect 3051 -1204 3085 -1188
rect 3169 1188 3203 1204
rect 3169 -1204 3203 -1188
rect 3287 1188 3321 1204
rect 3287 -1204 3321 -1188
rect 3405 1188 3439 1204
rect 3405 -1204 3439 -1188
rect 3523 1188 3557 1204
rect 3523 -1204 3557 -1188
rect 3641 1188 3675 1204
rect 3641 -1204 3675 -1188
rect 3759 1188 3793 1204
rect 3759 -1204 3793 -1188
rect 3877 1188 3911 1204
rect 3877 -1204 3911 -1188
rect 3995 1188 4029 1204
rect 3995 -1204 4029 -1188
rect 4113 1188 4147 1204
rect 4113 -1204 4147 -1188
rect 4231 1188 4265 1204
rect 4231 -1204 4265 -1188
rect 4349 1188 4383 1204
rect 4349 -1204 4383 -1188
rect 4467 1188 4501 1204
rect 4467 -1204 4501 -1188
rect 4585 1188 4619 1204
rect 4585 -1204 4619 -1188
rect 4703 1188 4737 1204
rect 4703 -1204 4737 -1188
rect 4821 1188 4855 1204
rect 4821 -1204 4855 -1188
rect 4939 1188 4973 1204
rect 4939 -1204 4973 -1188
rect 5057 1188 5091 1204
rect 5057 -1204 5091 -1188
rect 5175 1188 5209 1204
rect 5175 -1204 5209 -1188
rect 5293 1188 5327 1204
rect 5293 -1204 5327 -1188
rect -5284 -1272 -5268 -1238
rect -5234 -1272 -5218 -1238
rect -5166 -1272 -5150 -1238
rect -5116 -1272 -5100 -1238
rect -5048 -1272 -5032 -1238
rect -4998 -1272 -4982 -1238
rect -4930 -1272 -4914 -1238
rect -4880 -1272 -4864 -1238
rect -4812 -1272 -4796 -1238
rect -4762 -1272 -4746 -1238
rect -4694 -1272 -4678 -1238
rect -4644 -1272 -4628 -1238
rect -4576 -1272 -4560 -1238
rect -4526 -1272 -4510 -1238
rect -4458 -1272 -4442 -1238
rect -4408 -1272 -4392 -1238
rect -4340 -1272 -4324 -1238
rect -4290 -1272 -4274 -1238
rect -4222 -1272 -4206 -1238
rect -4172 -1272 -4156 -1238
rect -4104 -1272 -4088 -1238
rect -4054 -1272 -4038 -1238
rect -3986 -1272 -3970 -1238
rect -3936 -1272 -3920 -1238
rect -3868 -1272 -3852 -1238
rect -3818 -1272 -3802 -1238
rect -3750 -1272 -3734 -1238
rect -3700 -1272 -3684 -1238
rect -3632 -1272 -3616 -1238
rect -3582 -1272 -3566 -1238
rect -3514 -1272 -3498 -1238
rect -3464 -1272 -3448 -1238
rect -3396 -1272 -3380 -1238
rect -3346 -1272 -3330 -1238
rect -3278 -1272 -3262 -1238
rect -3228 -1272 -3212 -1238
rect -3160 -1272 -3144 -1238
rect -3110 -1272 -3094 -1238
rect -3042 -1272 -3026 -1238
rect -2992 -1272 -2976 -1238
rect -2924 -1272 -2908 -1238
rect -2874 -1272 -2858 -1238
rect -2806 -1272 -2790 -1238
rect -2756 -1272 -2740 -1238
rect -2688 -1272 -2672 -1238
rect -2638 -1272 -2622 -1238
rect -2570 -1272 -2554 -1238
rect -2520 -1272 -2504 -1238
rect -2452 -1272 -2436 -1238
rect -2402 -1272 -2386 -1238
rect -2334 -1272 -2318 -1238
rect -2284 -1272 -2268 -1238
rect -2216 -1272 -2200 -1238
rect -2166 -1272 -2150 -1238
rect -2098 -1272 -2082 -1238
rect -2048 -1272 -2032 -1238
rect -1980 -1272 -1964 -1238
rect -1930 -1272 -1914 -1238
rect -1862 -1272 -1846 -1238
rect -1812 -1272 -1796 -1238
rect -1744 -1272 -1728 -1238
rect -1694 -1272 -1678 -1238
rect -1626 -1272 -1610 -1238
rect -1576 -1272 -1560 -1238
rect -1508 -1272 -1492 -1238
rect -1458 -1272 -1442 -1238
rect -1390 -1272 -1374 -1238
rect -1340 -1272 -1324 -1238
rect -1272 -1272 -1256 -1238
rect -1222 -1272 -1206 -1238
rect -1154 -1272 -1138 -1238
rect -1104 -1272 -1088 -1238
rect -1036 -1272 -1020 -1238
rect -986 -1272 -970 -1238
rect -918 -1272 -902 -1238
rect -868 -1272 -852 -1238
rect -800 -1272 -784 -1238
rect -750 -1272 -734 -1238
rect -682 -1272 -666 -1238
rect -632 -1272 -616 -1238
rect -564 -1272 -548 -1238
rect -514 -1272 -498 -1238
rect -446 -1272 -430 -1238
rect -396 -1272 -380 -1238
rect -328 -1272 -312 -1238
rect -278 -1272 -262 -1238
rect -210 -1272 -194 -1238
rect -160 -1272 -144 -1238
rect -92 -1272 -76 -1238
rect -42 -1272 -26 -1238
rect 26 -1272 42 -1238
rect 76 -1272 92 -1238
rect 144 -1272 160 -1238
rect 194 -1272 210 -1238
rect 262 -1272 278 -1238
rect 312 -1272 328 -1238
rect 380 -1272 396 -1238
rect 430 -1272 446 -1238
rect 498 -1272 514 -1238
rect 548 -1272 564 -1238
rect 616 -1272 632 -1238
rect 666 -1272 682 -1238
rect 734 -1272 750 -1238
rect 784 -1272 800 -1238
rect 852 -1272 868 -1238
rect 902 -1272 918 -1238
rect 970 -1272 986 -1238
rect 1020 -1272 1036 -1238
rect 1088 -1272 1104 -1238
rect 1138 -1272 1154 -1238
rect 1206 -1272 1222 -1238
rect 1256 -1272 1272 -1238
rect 1324 -1272 1340 -1238
rect 1374 -1272 1390 -1238
rect 1442 -1272 1458 -1238
rect 1492 -1272 1508 -1238
rect 1560 -1272 1576 -1238
rect 1610 -1272 1626 -1238
rect 1678 -1272 1694 -1238
rect 1728 -1272 1744 -1238
rect 1796 -1272 1812 -1238
rect 1846 -1272 1862 -1238
rect 1914 -1272 1930 -1238
rect 1964 -1272 1980 -1238
rect 2032 -1272 2048 -1238
rect 2082 -1272 2098 -1238
rect 2150 -1272 2166 -1238
rect 2200 -1272 2216 -1238
rect 2268 -1272 2284 -1238
rect 2318 -1272 2334 -1238
rect 2386 -1272 2402 -1238
rect 2436 -1272 2452 -1238
rect 2504 -1272 2520 -1238
rect 2554 -1272 2570 -1238
rect 2622 -1272 2638 -1238
rect 2672 -1272 2688 -1238
rect 2740 -1272 2756 -1238
rect 2790 -1272 2806 -1238
rect 2858 -1272 2874 -1238
rect 2908 -1272 2924 -1238
rect 2976 -1272 2992 -1238
rect 3026 -1272 3042 -1238
rect 3094 -1272 3110 -1238
rect 3144 -1272 3160 -1238
rect 3212 -1272 3228 -1238
rect 3262 -1272 3278 -1238
rect 3330 -1272 3346 -1238
rect 3380 -1272 3396 -1238
rect 3448 -1272 3464 -1238
rect 3498 -1272 3514 -1238
rect 3566 -1272 3582 -1238
rect 3616 -1272 3632 -1238
rect 3684 -1272 3700 -1238
rect 3734 -1272 3750 -1238
rect 3802 -1272 3818 -1238
rect 3852 -1272 3868 -1238
rect 3920 -1272 3936 -1238
rect 3970 -1272 3986 -1238
rect 4038 -1272 4054 -1238
rect 4088 -1272 4104 -1238
rect 4156 -1272 4172 -1238
rect 4206 -1272 4222 -1238
rect 4274 -1272 4290 -1238
rect 4324 -1272 4340 -1238
rect 4392 -1272 4408 -1238
rect 4442 -1272 4458 -1238
rect 4510 -1272 4526 -1238
rect 4560 -1272 4576 -1238
rect 4628 -1272 4644 -1238
rect 4678 -1272 4694 -1238
rect 4746 -1272 4762 -1238
rect 4796 -1272 4812 -1238
rect 4864 -1272 4880 -1238
rect 4914 -1272 4930 -1238
rect 4982 -1272 4998 -1238
rect 5032 -1272 5048 -1238
rect 5100 -1272 5116 -1238
rect 5150 -1272 5166 -1238
rect 5218 -1272 5234 -1238
rect 5268 -1272 5284 -1238
rect -5441 -1340 -5407 -1278
rect 5407 -1340 5441 -1278
rect -5441 -1374 -5345 -1340
rect 5345 -1374 5441 -1340
<< viali >>
rect -5268 1238 -5234 1272
rect -5150 1238 -5116 1272
rect -5032 1238 -4998 1272
rect -4914 1238 -4880 1272
rect -4796 1238 -4762 1272
rect -4678 1238 -4644 1272
rect -4560 1238 -4526 1272
rect -4442 1238 -4408 1272
rect -4324 1238 -4290 1272
rect -4206 1238 -4172 1272
rect -4088 1238 -4054 1272
rect -3970 1238 -3936 1272
rect -3852 1238 -3818 1272
rect -3734 1238 -3700 1272
rect -3616 1238 -3582 1272
rect -3498 1238 -3464 1272
rect -3380 1238 -3346 1272
rect -3262 1238 -3228 1272
rect -3144 1238 -3110 1272
rect -3026 1238 -2992 1272
rect -2908 1238 -2874 1272
rect -2790 1238 -2756 1272
rect -2672 1238 -2638 1272
rect -2554 1238 -2520 1272
rect -2436 1238 -2402 1272
rect -2318 1238 -2284 1272
rect -2200 1238 -2166 1272
rect -2082 1238 -2048 1272
rect -1964 1238 -1930 1272
rect -1846 1238 -1812 1272
rect -1728 1238 -1694 1272
rect -1610 1238 -1576 1272
rect -1492 1238 -1458 1272
rect -1374 1238 -1340 1272
rect -1256 1238 -1222 1272
rect -1138 1238 -1104 1272
rect -1020 1238 -986 1272
rect -902 1238 -868 1272
rect -784 1238 -750 1272
rect -666 1238 -632 1272
rect -548 1238 -514 1272
rect -430 1238 -396 1272
rect -312 1238 -278 1272
rect -194 1238 -160 1272
rect -76 1238 -42 1272
rect 42 1238 76 1272
rect 160 1238 194 1272
rect 278 1238 312 1272
rect 396 1238 430 1272
rect 514 1238 548 1272
rect 632 1238 666 1272
rect 750 1238 784 1272
rect 868 1238 902 1272
rect 986 1238 1020 1272
rect 1104 1238 1138 1272
rect 1222 1238 1256 1272
rect 1340 1238 1374 1272
rect 1458 1238 1492 1272
rect 1576 1238 1610 1272
rect 1694 1238 1728 1272
rect 1812 1238 1846 1272
rect 1930 1238 1964 1272
rect 2048 1238 2082 1272
rect 2166 1238 2200 1272
rect 2284 1238 2318 1272
rect 2402 1238 2436 1272
rect 2520 1238 2554 1272
rect 2638 1238 2672 1272
rect 2756 1238 2790 1272
rect 2874 1238 2908 1272
rect 2992 1238 3026 1272
rect 3110 1238 3144 1272
rect 3228 1238 3262 1272
rect 3346 1238 3380 1272
rect 3464 1238 3498 1272
rect 3582 1238 3616 1272
rect 3700 1238 3734 1272
rect 3818 1238 3852 1272
rect 3936 1238 3970 1272
rect 4054 1238 4088 1272
rect 4172 1238 4206 1272
rect 4290 1238 4324 1272
rect 4408 1238 4442 1272
rect 4526 1238 4560 1272
rect 4644 1238 4678 1272
rect 4762 1238 4796 1272
rect 4880 1238 4914 1272
rect 4998 1238 5032 1272
rect 5116 1238 5150 1272
rect 5234 1238 5268 1272
rect -5327 -1188 -5293 1188
rect -5209 -1188 -5175 1188
rect -5091 -1188 -5057 1188
rect -4973 -1188 -4939 1188
rect -4855 -1188 -4821 1188
rect -4737 -1188 -4703 1188
rect -4619 -1188 -4585 1188
rect -4501 -1188 -4467 1188
rect -4383 -1188 -4349 1188
rect -4265 -1188 -4231 1188
rect -4147 -1188 -4113 1188
rect -4029 -1188 -3995 1188
rect -3911 -1188 -3877 1188
rect -3793 -1188 -3759 1188
rect -3675 -1188 -3641 1188
rect -3557 -1188 -3523 1188
rect -3439 -1188 -3405 1188
rect -3321 -1188 -3287 1188
rect -3203 -1188 -3169 1188
rect -3085 -1188 -3051 1188
rect -2967 -1188 -2933 1188
rect -2849 -1188 -2815 1188
rect -2731 -1188 -2697 1188
rect -2613 -1188 -2579 1188
rect -2495 -1188 -2461 1188
rect -2377 -1188 -2343 1188
rect -2259 -1188 -2225 1188
rect -2141 -1188 -2107 1188
rect -2023 -1188 -1989 1188
rect -1905 -1188 -1871 1188
rect -1787 -1188 -1753 1188
rect -1669 -1188 -1635 1188
rect -1551 -1188 -1517 1188
rect -1433 -1188 -1399 1188
rect -1315 -1188 -1281 1188
rect -1197 -1188 -1163 1188
rect -1079 -1188 -1045 1188
rect -961 -1188 -927 1188
rect -843 -1188 -809 1188
rect -725 -1188 -691 1188
rect -607 -1188 -573 1188
rect -489 -1188 -455 1188
rect -371 -1188 -337 1188
rect -253 -1188 -219 1188
rect -135 -1188 -101 1188
rect -17 -1188 17 1188
rect 101 -1188 135 1188
rect 219 -1188 253 1188
rect 337 -1188 371 1188
rect 455 -1188 489 1188
rect 573 -1188 607 1188
rect 691 -1188 725 1188
rect 809 -1188 843 1188
rect 927 -1188 961 1188
rect 1045 -1188 1079 1188
rect 1163 -1188 1197 1188
rect 1281 -1188 1315 1188
rect 1399 -1188 1433 1188
rect 1517 -1188 1551 1188
rect 1635 -1188 1669 1188
rect 1753 -1188 1787 1188
rect 1871 -1188 1905 1188
rect 1989 -1188 2023 1188
rect 2107 -1188 2141 1188
rect 2225 -1188 2259 1188
rect 2343 -1188 2377 1188
rect 2461 -1188 2495 1188
rect 2579 -1188 2613 1188
rect 2697 -1188 2731 1188
rect 2815 -1188 2849 1188
rect 2933 -1188 2967 1188
rect 3051 -1188 3085 1188
rect 3169 -1188 3203 1188
rect 3287 -1188 3321 1188
rect 3405 -1188 3439 1188
rect 3523 -1188 3557 1188
rect 3641 -1188 3675 1188
rect 3759 -1188 3793 1188
rect 3877 -1188 3911 1188
rect 3995 -1188 4029 1188
rect 4113 -1188 4147 1188
rect 4231 -1188 4265 1188
rect 4349 -1188 4383 1188
rect 4467 -1188 4501 1188
rect 4585 -1188 4619 1188
rect 4703 -1188 4737 1188
rect 4821 -1188 4855 1188
rect 4939 -1188 4973 1188
rect 5057 -1188 5091 1188
rect 5175 -1188 5209 1188
rect 5293 -1188 5327 1188
rect -5268 -1272 -5234 -1238
rect -5150 -1272 -5116 -1238
rect -5032 -1272 -4998 -1238
rect -4914 -1272 -4880 -1238
rect -4796 -1272 -4762 -1238
rect -4678 -1272 -4644 -1238
rect -4560 -1272 -4526 -1238
rect -4442 -1272 -4408 -1238
rect -4324 -1272 -4290 -1238
rect -4206 -1272 -4172 -1238
rect -4088 -1272 -4054 -1238
rect -3970 -1272 -3936 -1238
rect -3852 -1272 -3818 -1238
rect -3734 -1272 -3700 -1238
rect -3616 -1272 -3582 -1238
rect -3498 -1272 -3464 -1238
rect -3380 -1272 -3346 -1238
rect -3262 -1272 -3228 -1238
rect -3144 -1272 -3110 -1238
rect -3026 -1272 -2992 -1238
rect -2908 -1272 -2874 -1238
rect -2790 -1272 -2756 -1238
rect -2672 -1272 -2638 -1238
rect -2554 -1272 -2520 -1238
rect -2436 -1272 -2402 -1238
rect -2318 -1272 -2284 -1238
rect -2200 -1272 -2166 -1238
rect -2082 -1272 -2048 -1238
rect -1964 -1272 -1930 -1238
rect -1846 -1272 -1812 -1238
rect -1728 -1272 -1694 -1238
rect -1610 -1272 -1576 -1238
rect -1492 -1272 -1458 -1238
rect -1374 -1272 -1340 -1238
rect -1256 -1272 -1222 -1238
rect -1138 -1272 -1104 -1238
rect -1020 -1272 -986 -1238
rect -902 -1272 -868 -1238
rect -784 -1272 -750 -1238
rect -666 -1272 -632 -1238
rect -548 -1272 -514 -1238
rect -430 -1272 -396 -1238
rect -312 -1272 -278 -1238
rect -194 -1272 -160 -1238
rect -76 -1272 -42 -1238
rect 42 -1272 76 -1238
rect 160 -1272 194 -1238
rect 278 -1272 312 -1238
rect 396 -1272 430 -1238
rect 514 -1272 548 -1238
rect 632 -1272 666 -1238
rect 750 -1272 784 -1238
rect 868 -1272 902 -1238
rect 986 -1272 1020 -1238
rect 1104 -1272 1138 -1238
rect 1222 -1272 1256 -1238
rect 1340 -1272 1374 -1238
rect 1458 -1272 1492 -1238
rect 1576 -1272 1610 -1238
rect 1694 -1272 1728 -1238
rect 1812 -1272 1846 -1238
rect 1930 -1272 1964 -1238
rect 2048 -1272 2082 -1238
rect 2166 -1272 2200 -1238
rect 2284 -1272 2318 -1238
rect 2402 -1272 2436 -1238
rect 2520 -1272 2554 -1238
rect 2638 -1272 2672 -1238
rect 2756 -1272 2790 -1238
rect 2874 -1272 2908 -1238
rect 2992 -1272 3026 -1238
rect 3110 -1272 3144 -1238
rect 3228 -1272 3262 -1238
rect 3346 -1272 3380 -1238
rect 3464 -1272 3498 -1238
rect 3582 -1272 3616 -1238
rect 3700 -1272 3734 -1238
rect 3818 -1272 3852 -1238
rect 3936 -1272 3970 -1238
rect 4054 -1272 4088 -1238
rect 4172 -1272 4206 -1238
rect 4290 -1272 4324 -1238
rect 4408 -1272 4442 -1238
rect 4526 -1272 4560 -1238
rect 4644 -1272 4678 -1238
rect 4762 -1272 4796 -1238
rect 4880 -1272 4914 -1238
rect 4998 -1272 5032 -1238
rect 5116 -1272 5150 -1238
rect 5234 -1272 5268 -1238
<< metal1 >>
rect -5280 1272 -5222 1278
rect -5280 1238 -5268 1272
rect -5234 1238 -5222 1272
rect -5280 1232 -5222 1238
rect -5162 1272 -5104 1278
rect -5162 1238 -5150 1272
rect -5116 1238 -5104 1272
rect -5162 1232 -5104 1238
rect -5044 1272 -4986 1278
rect -5044 1238 -5032 1272
rect -4998 1238 -4986 1272
rect -5044 1232 -4986 1238
rect -4926 1272 -4868 1278
rect -4926 1238 -4914 1272
rect -4880 1238 -4868 1272
rect -4926 1232 -4868 1238
rect -4808 1272 -4750 1278
rect -4808 1238 -4796 1272
rect -4762 1238 -4750 1272
rect -4808 1232 -4750 1238
rect -4690 1272 -4632 1278
rect -4690 1238 -4678 1272
rect -4644 1238 -4632 1272
rect -4690 1232 -4632 1238
rect -4572 1272 -4514 1278
rect -4572 1238 -4560 1272
rect -4526 1238 -4514 1272
rect -4572 1232 -4514 1238
rect -4454 1272 -4396 1278
rect -4454 1238 -4442 1272
rect -4408 1238 -4396 1272
rect -4454 1232 -4396 1238
rect -4336 1272 -4278 1278
rect -4336 1238 -4324 1272
rect -4290 1238 -4278 1272
rect -4336 1232 -4278 1238
rect -4218 1272 -4160 1278
rect -4218 1238 -4206 1272
rect -4172 1238 -4160 1272
rect -4218 1232 -4160 1238
rect -4100 1272 -4042 1278
rect -4100 1238 -4088 1272
rect -4054 1238 -4042 1272
rect -4100 1232 -4042 1238
rect -3982 1272 -3924 1278
rect -3982 1238 -3970 1272
rect -3936 1238 -3924 1272
rect -3982 1232 -3924 1238
rect -3864 1272 -3806 1278
rect -3864 1238 -3852 1272
rect -3818 1238 -3806 1272
rect -3864 1232 -3806 1238
rect -3746 1272 -3688 1278
rect -3746 1238 -3734 1272
rect -3700 1238 -3688 1272
rect -3746 1232 -3688 1238
rect -3628 1272 -3570 1278
rect -3628 1238 -3616 1272
rect -3582 1238 -3570 1272
rect -3628 1232 -3570 1238
rect -3510 1272 -3452 1278
rect -3510 1238 -3498 1272
rect -3464 1238 -3452 1272
rect -3510 1232 -3452 1238
rect -3392 1272 -3334 1278
rect -3392 1238 -3380 1272
rect -3346 1238 -3334 1272
rect -3392 1232 -3334 1238
rect -3274 1272 -3216 1278
rect -3274 1238 -3262 1272
rect -3228 1238 -3216 1272
rect -3274 1232 -3216 1238
rect -3156 1272 -3098 1278
rect -3156 1238 -3144 1272
rect -3110 1238 -3098 1272
rect -3156 1232 -3098 1238
rect -3038 1272 -2980 1278
rect -3038 1238 -3026 1272
rect -2992 1238 -2980 1272
rect -3038 1232 -2980 1238
rect -2920 1272 -2862 1278
rect -2920 1238 -2908 1272
rect -2874 1238 -2862 1272
rect -2920 1232 -2862 1238
rect -2802 1272 -2744 1278
rect -2802 1238 -2790 1272
rect -2756 1238 -2744 1272
rect -2802 1232 -2744 1238
rect -2684 1272 -2626 1278
rect -2684 1238 -2672 1272
rect -2638 1238 -2626 1272
rect -2684 1232 -2626 1238
rect -2566 1272 -2508 1278
rect -2566 1238 -2554 1272
rect -2520 1238 -2508 1272
rect -2566 1232 -2508 1238
rect -2448 1272 -2390 1278
rect -2448 1238 -2436 1272
rect -2402 1238 -2390 1272
rect -2448 1232 -2390 1238
rect -2330 1272 -2272 1278
rect -2330 1238 -2318 1272
rect -2284 1238 -2272 1272
rect -2330 1232 -2272 1238
rect -2212 1272 -2154 1278
rect -2212 1238 -2200 1272
rect -2166 1238 -2154 1272
rect -2212 1232 -2154 1238
rect -2094 1272 -2036 1278
rect -2094 1238 -2082 1272
rect -2048 1238 -2036 1272
rect -2094 1232 -2036 1238
rect -1976 1272 -1918 1278
rect -1976 1238 -1964 1272
rect -1930 1238 -1918 1272
rect -1976 1232 -1918 1238
rect -1858 1272 -1800 1278
rect -1858 1238 -1846 1272
rect -1812 1238 -1800 1272
rect -1858 1232 -1800 1238
rect -1740 1272 -1682 1278
rect -1740 1238 -1728 1272
rect -1694 1238 -1682 1272
rect -1740 1232 -1682 1238
rect -1622 1272 -1564 1278
rect -1622 1238 -1610 1272
rect -1576 1238 -1564 1272
rect -1622 1232 -1564 1238
rect -1504 1272 -1446 1278
rect -1504 1238 -1492 1272
rect -1458 1238 -1446 1272
rect -1504 1232 -1446 1238
rect -1386 1272 -1328 1278
rect -1386 1238 -1374 1272
rect -1340 1238 -1328 1272
rect -1386 1232 -1328 1238
rect -1268 1272 -1210 1278
rect -1268 1238 -1256 1272
rect -1222 1238 -1210 1272
rect -1268 1232 -1210 1238
rect -1150 1272 -1092 1278
rect -1150 1238 -1138 1272
rect -1104 1238 -1092 1272
rect -1150 1232 -1092 1238
rect -1032 1272 -974 1278
rect -1032 1238 -1020 1272
rect -986 1238 -974 1272
rect -1032 1232 -974 1238
rect -914 1272 -856 1278
rect -914 1238 -902 1272
rect -868 1238 -856 1272
rect -914 1232 -856 1238
rect -796 1272 -738 1278
rect -796 1238 -784 1272
rect -750 1238 -738 1272
rect -796 1232 -738 1238
rect -678 1272 -620 1278
rect -678 1238 -666 1272
rect -632 1238 -620 1272
rect -678 1232 -620 1238
rect -560 1272 -502 1278
rect -560 1238 -548 1272
rect -514 1238 -502 1272
rect -560 1232 -502 1238
rect -442 1272 -384 1278
rect -442 1238 -430 1272
rect -396 1238 -384 1272
rect -442 1232 -384 1238
rect -324 1272 -266 1278
rect -324 1238 -312 1272
rect -278 1238 -266 1272
rect -324 1232 -266 1238
rect -206 1272 -148 1278
rect -206 1238 -194 1272
rect -160 1238 -148 1272
rect -206 1232 -148 1238
rect -88 1272 -30 1278
rect -88 1238 -76 1272
rect -42 1238 -30 1272
rect -88 1232 -30 1238
rect 30 1272 88 1278
rect 30 1238 42 1272
rect 76 1238 88 1272
rect 30 1232 88 1238
rect 148 1272 206 1278
rect 148 1238 160 1272
rect 194 1238 206 1272
rect 148 1232 206 1238
rect 266 1272 324 1278
rect 266 1238 278 1272
rect 312 1238 324 1272
rect 266 1232 324 1238
rect 384 1272 442 1278
rect 384 1238 396 1272
rect 430 1238 442 1272
rect 384 1232 442 1238
rect 502 1272 560 1278
rect 502 1238 514 1272
rect 548 1238 560 1272
rect 502 1232 560 1238
rect 620 1272 678 1278
rect 620 1238 632 1272
rect 666 1238 678 1272
rect 620 1232 678 1238
rect 738 1272 796 1278
rect 738 1238 750 1272
rect 784 1238 796 1272
rect 738 1232 796 1238
rect 856 1272 914 1278
rect 856 1238 868 1272
rect 902 1238 914 1272
rect 856 1232 914 1238
rect 974 1272 1032 1278
rect 974 1238 986 1272
rect 1020 1238 1032 1272
rect 974 1232 1032 1238
rect 1092 1272 1150 1278
rect 1092 1238 1104 1272
rect 1138 1238 1150 1272
rect 1092 1232 1150 1238
rect 1210 1272 1268 1278
rect 1210 1238 1222 1272
rect 1256 1238 1268 1272
rect 1210 1232 1268 1238
rect 1328 1272 1386 1278
rect 1328 1238 1340 1272
rect 1374 1238 1386 1272
rect 1328 1232 1386 1238
rect 1446 1272 1504 1278
rect 1446 1238 1458 1272
rect 1492 1238 1504 1272
rect 1446 1232 1504 1238
rect 1564 1272 1622 1278
rect 1564 1238 1576 1272
rect 1610 1238 1622 1272
rect 1564 1232 1622 1238
rect 1682 1272 1740 1278
rect 1682 1238 1694 1272
rect 1728 1238 1740 1272
rect 1682 1232 1740 1238
rect 1800 1272 1858 1278
rect 1800 1238 1812 1272
rect 1846 1238 1858 1272
rect 1800 1232 1858 1238
rect 1918 1272 1976 1278
rect 1918 1238 1930 1272
rect 1964 1238 1976 1272
rect 1918 1232 1976 1238
rect 2036 1272 2094 1278
rect 2036 1238 2048 1272
rect 2082 1238 2094 1272
rect 2036 1232 2094 1238
rect 2154 1272 2212 1278
rect 2154 1238 2166 1272
rect 2200 1238 2212 1272
rect 2154 1232 2212 1238
rect 2272 1272 2330 1278
rect 2272 1238 2284 1272
rect 2318 1238 2330 1272
rect 2272 1232 2330 1238
rect 2390 1272 2448 1278
rect 2390 1238 2402 1272
rect 2436 1238 2448 1272
rect 2390 1232 2448 1238
rect 2508 1272 2566 1278
rect 2508 1238 2520 1272
rect 2554 1238 2566 1272
rect 2508 1232 2566 1238
rect 2626 1272 2684 1278
rect 2626 1238 2638 1272
rect 2672 1238 2684 1272
rect 2626 1232 2684 1238
rect 2744 1272 2802 1278
rect 2744 1238 2756 1272
rect 2790 1238 2802 1272
rect 2744 1232 2802 1238
rect 2862 1272 2920 1278
rect 2862 1238 2874 1272
rect 2908 1238 2920 1272
rect 2862 1232 2920 1238
rect 2980 1272 3038 1278
rect 2980 1238 2992 1272
rect 3026 1238 3038 1272
rect 2980 1232 3038 1238
rect 3098 1272 3156 1278
rect 3098 1238 3110 1272
rect 3144 1238 3156 1272
rect 3098 1232 3156 1238
rect 3216 1272 3274 1278
rect 3216 1238 3228 1272
rect 3262 1238 3274 1272
rect 3216 1232 3274 1238
rect 3334 1272 3392 1278
rect 3334 1238 3346 1272
rect 3380 1238 3392 1272
rect 3334 1232 3392 1238
rect 3452 1272 3510 1278
rect 3452 1238 3464 1272
rect 3498 1238 3510 1272
rect 3452 1232 3510 1238
rect 3570 1272 3628 1278
rect 3570 1238 3582 1272
rect 3616 1238 3628 1272
rect 3570 1232 3628 1238
rect 3688 1272 3746 1278
rect 3688 1238 3700 1272
rect 3734 1238 3746 1272
rect 3688 1232 3746 1238
rect 3806 1272 3864 1278
rect 3806 1238 3818 1272
rect 3852 1238 3864 1272
rect 3806 1232 3864 1238
rect 3924 1272 3982 1278
rect 3924 1238 3936 1272
rect 3970 1238 3982 1272
rect 3924 1232 3982 1238
rect 4042 1272 4100 1278
rect 4042 1238 4054 1272
rect 4088 1238 4100 1272
rect 4042 1232 4100 1238
rect 4160 1272 4218 1278
rect 4160 1238 4172 1272
rect 4206 1238 4218 1272
rect 4160 1232 4218 1238
rect 4278 1272 4336 1278
rect 4278 1238 4290 1272
rect 4324 1238 4336 1272
rect 4278 1232 4336 1238
rect 4396 1272 4454 1278
rect 4396 1238 4408 1272
rect 4442 1238 4454 1272
rect 4396 1232 4454 1238
rect 4514 1272 4572 1278
rect 4514 1238 4526 1272
rect 4560 1238 4572 1272
rect 4514 1232 4572 1238
rect 4632 1272 4690 1278
rect 4632 1238 4644 1272
rect 4678 1238 4690 1272
rect 4632 1232 4690 1238
rect 4750 1272 4808 1278
rect 4750 1238 4762 1272
rect 4796 1238 4808 1272
rect 4750 1232 4808 1238
rect 4868 1272 4926 1278
rect 4868 1238 4880 1272
rect 4914 1238 4926 1272
rect 4868 1232 4926 1238
rect 4986 1272 5044 1278
rect 4986 1238 4998 1272
rect 5032 1238 5044 1272
rect 4986 1232 5044 1238
rect 5104 1272 5162 1278
rect 5104 1238 5116 1272
rect 5150 1238 5162 1272
rect 5104 1232 5162 1238
rect 5222 1272 5280 1278
rect 5222 1238 5234 1272
rect 5268 1238 5280 1272
rect 5222 1232 5280 1238
rect -5333 1188 -5287 1200
rect -5333 -1188 -5327 1188
rect -5293 -1188 -5287 1188
rect -5333 -1200 -5287 -1188
rect -5215 1188 -5169 1200
rect -5215 -1188 -5209 1188
rect -5175 -1188 -5169 1188
rect -5215 -1200 -5169 -1188
rect -5097 1188 -5051 1200
rect -5097 -1188 -5091 1188
rect -5057 -1188 -5051 1188
rect -5097 -1200 -5051 -1188
rect -4979 1188 -4933 1200
rect -4979 -1188 -4973 1188
rect -4939 -1188 -4933 1188
rect -4979 -1200 -4933 -1188
rect -4861 1188 -4815 1200
rect -4861 -1188 -4855 1188
rect -4821 -1188 -4815 1188
rect -4861 -1200 -4815 -1188
rect -4743 1188 -4697 1200
rect -4743 -1188 -4737 1188
rect -4703 -1188 -4697 1188
rect -4743 -1200 -4697 -1188
rect -4625 1188 -4579 1200
rect -4625 -1188 -4619 1188
rect -4585 -1188 -4579 1188
rect -4625 -1200 -4579 -1188
rect -4507 1188 -4461 1200
rect -4507 -1188 -4501 1188
rect -4467 -1188 -4461 1188
rect -4507 -1200 -4461 -1188
rect -4389 1188 -4343 1200
rect -4389 -1188 -4383 1188
rect -4349 -1188 -4343 1188
rect -4389 -1200 -4343 -1188
rect -4271 1188 -4225 1200
rect -4271 -1188 -4265 1188
rect -4231 -1188 -4225 1188
rect -4271 -1200 -4225 -1188
rect -4153 1188 -4107 1200
rect -4153 -1188 -4147 1188
rect -4113 -1188 -4107 1188
rect -4153 -1200 -4107 -1188
rect -4035 1188 -3989 1200
rect -4035 -1188 -4029 1188
rect -3995 -1188 -3989 1188
rect -4035 -1200 -3989 -1188
rect -3917 1188 -3871 1200
rect -3917 -1188 -3911 1188
rect -3877 -1188 -3871 1188
rect -3917 -1200 -3871 -1188
rect -3799 1188 -3753 1200
rect -3799 -1188 -3793 1188
rect -3759 -1188 -3753 1188
rect -3799 -1200 -3753 -1188
rect -3681 1188 -3635 1200
rect -3681 -1188 -3675 1188
rect -3641 -1188 -3635 1188
rect -3681 -1200 -3635 -1188
rect -3563 1188 -3517 1200
rect -3563 -1188 -3557 1188
rect -3523 -1188 -3517 1188
rect -3563 -1200 -3517 -1188
rect -3445 1188 -3399 1200
rect -3445 -1188 -3439 1188
rect -3405 -1188 -3399 1188
rect -3445 -1200 -3399 -1188
rect -3327 1188 -3281 1200
rect -3327 -1188 -3321 1188
rect -3287 -1188 -3281 1188
rect -3327 -1200 -3281 -1188
rect -3209 1188 -3163 1200
rect -3209 -1188 -3203 1188
rect -3169 -1188 -3163 1188
rect -3209 -1200 -3163 -1188
rect -3091 1188 -3045 1200
rect -3091 -1188 -3085 1188
rect -3051 -1188 -3045 1188
rect -3091 -1200 -3045 -1188
rect -2973 1188 -2927 1200
rect -2973 -1188 -2967 1188
rect -2933 -1188 -2927 1188
rect -2973 -1200 -2927 -1188
rect -2855 1188 -2809 1200
rect -2855 -1188 -2849 1188
rect -2815 -1188 -2809 1188
rect -2855 -1200 -2809 -1188
rect -2737 1188 -2691 1200
rect -2737 -1188 -2731 1188
rect -2697 -1188 -2691 1188
rect -2737 -1200 -2691 -1188
rect -2619 1188 -2573 1200
rect -2619 -1188 -2613 1188
rect -2579 -1188 -2573 1188
rect -2619 -1200 -2573 -1188
rect -2501 1188 -2455 1200
rect -2501 -1188 -2495 1188
rect -2461 -1188 -2455 1188
rect -2501 -1200 -2455 -1188
rect -2383 1188 -2337 1200
rect -2383 -1188 -2377 1188
rect -2343 -1188 -2337 1188
rect -2383 -1200 -2337 -1188
rect -2265 1188 -2219 1200
rect -2265 -1188 -2259 1188
rect -2225 -1188 -2219 1188
rect -2265 -1200 -2219 -1188
rect -2147 1188 -2101 1200
rect -2147 -1188 -2141 1188
rect -2107 -1188 -2101 1188
rect -2147 -1200 -2101 -1188
rect -2029 1188 -1983 1200
rect -2029 -1188 -2023 1188
rect -1989 -1188 -1983 1188
rect -2029 -1200 -1983 -1188
rect -1911 1188 -1865 1200
rect -1911 -1188 -1905 1188
rect -1871 -1188 -1865 1188
rect -1911 -1200 -1865 -1188
rect -1793 1188 -1747 1200
rect -1793 -1188 -1787 1188
rect -1753 -1188 -1747 1188
rect -1793 -1200 -1747 -1188
rect -1675 1188 -1629 1200
rect -1675 -1188 -1669 1188
rect -1635 -1188 -1629 1188
rect -1675 -1200 -1629 -1188
rect -1557 1188 -1511 1200
rect -1557 -1188 -1551 1188
rect -1517 -1188 -1511 1188
rect -1557 -1200 -1511 -1188
rect -1439 1188 -1393 1200
rect -1439 -1188 -1433 1188
rect -1399 -1188 -1393 1188
rect -1439 -1200 -1393 -1188
rect -1321 1188 -1275 1200
rect -1321 -1188 -1315 1188
rect -1281 -1188 -1275 1188
rect -1321 -1200 -1275 -1188
rect -1203 1188 -1157 1200
rect -1203 -1188 -1197 1188
rect -1163 -1188 -1157 1188
rect -1203 -1200 -1157 -1188
rect -1085 1188 -1039 1200
rect -1085 -1188 -1079 1188
rect -1045 -1188 -1039 1188
rect -1085 -1200 -1039 -1188
rect -967 1188 -921 1200
rect -967 -1188 -961 1188
rect -927 -1188 -921 1188
rect -967 -1200 -921 -1188
rect -849 1188 -803 1200
rect -849 -1188 -843 1188
rect -809 -1188 -803 1188
rect -849 -1200 -803 -1188
rect -731 1188 -685 1200
rect -731 -1188 -725 1188
rect -691 -1188 -685 1188
rect -731 -1200 -685 -1188
rect -613 1188 -567 1200
rect -613 -1188 -607 1188
rect -573 -1188 -567 1188
rect -613 -1200 -567 -1188
rect -495 1188 -449 1200
rect -495 -1188 -489 1188
rect -455 -1188 -449 1188
rect -495 -1200 -449 -1188
rect -377 1188 -331 1200
rect -377 -1188 -371 1188
rect -337 -1188 -331 1188
rect -377 -1200 -331 -1188
rect -259 1188 -213 1200
rect -259 -1188 -253 1188
rect -219 -1188 -213 1188
rect -259 -1200 -213 -1188
rect -141 1188 -95 1200
rect -141 -1188 -135 1188
rect -101 -1188 -95 1188
rect -141 -1200 -95 -1188
rect -23 1188 23 1200
rect -23 -1188 -17 1188
rect 17 -1188 23 1188
rect -23 -1200 23 -1188
rect 95 1188 141 1200
rect 95 -1188 101 1188
rect 135 -1188 141 1188
rect 95 -1200 141 -1188
rect 213 1188 259 1200
rect 213 -1188 219 1188
rect 253 -1188 259 1188
rect 213 -1200 259 -1188
rect 331 1188 377 1200
rect 331 -1188 337 1188
rect 371 -1188 377 1188
rect 331 -1200 377 -1188
rect 449 1188 495 1200
rect 449 -1188 455 1188
rect 489 -1188 495 1188
rect 449 -1200 495 -1188
rect 567 1188 613 1200
rect 567 -1188 573 1188
rect 607 -1188 613 1188
rect 567 -1200 613 -1188
rect 685 1188 731 1200
rect 685 -1188 691 1188
rect 725 -1188 731 1188
rect 685 -1200 731 -1188
rect 803 1188 849 1200
rect 803 -1188 809 1188
rect 843 -1188 849 1188
rect 803 -1200 849 -1188
rect 921 1188 967 1200
rect 921 -1188 927 1188
rect 961 -1188 967 1188
rect 921 -1200 967 -1188
rect 1039 1188 1085 1200
rect 1039 -1188 1045 1188
rect 1079 -1188 1085 1188
rect 1039 -1200 1085 -1188
rect 1157 1188 1203 1200
rect 1157 -1188 1163 1188
rect 1197 -1188 1203 1188
rect 1157 -1200 1203 -1188
rect 1275 1188 1321 1200
rect 1275 -1188 1281 1188
rect 1315 -1188 1321 1188
rect 1275 -1200 1321 -1188
rect 1393 1188 1439 1200
rect 1393 -1188 1399 1188
rect 1433 -1188 1439 1188
rect 1393 -1200 1439 -1188
rect 1511 1188 1557 1200
rect 1511 -1188 1517 1188
rect 1551 -1188 1557 1188
rect 1511 -1200 1557 -1188
rect 1629 1188 1675 1200
rect 1629 -1188 1635 1188
rect 1669 -1188 1675 1188
rect 1629 -1200 1675 -1188
rect 1747 1188 1793 1200
rect 1747 -1188 1753 1188
rect 1787 -1188 1793 1188
rect 1747 -1200 1793 -1188
rect 1865 1188 1911 1200
rect 1865 -1188 1871 1188
rect 1905 -1188 1911 1188
rect 1865 -1200 1911 -1188
rect 1983 1188 2029 1200
rect 1983 -1188 1989 1188
rect 2023 -1188 2029 1188
rect 1983 -1200 2029 -1188
rect 2101 1188 2147 1200
rect 2101 -1188 2107 1188
rect 2141 -1188 2147 1188
rect 2101 -1200 2147 -1188
rect 2219 1188 2265 1200
rect 2219 -1188 2225 1188
rect 2259 -1188 2265 1188
rect 2219 -1200 2265 -1188
rect 2337 1188 2383 1200
rect 2337 -1188 2343 1188
rect 2377 -1188 2383 1188
rect 2337 -1200 2383 -1188
rect 2455 1188 2501 1200
rect 2455 -1188 2461 1188
rect 2495 -1188 2501 1188
rect 2455 -1200 2501 -1188
rect 2573 1188 2619 1200
rect 2573 -1188 2579 1188
rect 2613 -1188 2619 1188
rect 2573 -1200 2619 -1188
rect 2691 1188 2737 1200
rect 2691 -1188 2697 1188
rect 2731 -1188 2737 1188
rect 2691 -1200 2737 -1188
rect 2809 1188 2855 1200
rect 2809 -1188 2815 1188
rect 2849 -1188 2855 1188
rect 2809 -1200 2855 -1188
rect 2927 1188 2973 1200
rect 2927 -1188 2933 1188
rect 2967 -1188 2973 1188
rect 2927 -1200 2973 -1188
rect 3045 1188 3091 1200
rect 3045 -1188 3051 1188
rect 3085 -1188 3091 1188
rect 3045 -1200 3091 -1188
rect 3163 1188 3209 1200
rect 3163 -1188 3169 1188
rect 3203 -1188 3209 1188
rect 3163 -1200 3209 -1188
rect 3281 1188 3327 1200
rect 3281 -1188 3287 1188
rect 3321 -1188 3327 1188
rect 3281 -1200 3327 -1188
rect 3399 1188 3445 1200
rect 3399 -1188 3405 1188
rect 3439 -1188 3445 1188
rect 3399 -1200 3445 -1188
rect 3517 1188 3563 1200
rect 3517 -1188 3523 1188
rect 3557 -1188 3563 1188
rect 3517 -1200 3563 -1188
rect 3635 1188 3681 1200
rect 3635 -1188 3641 1188
rect 3675 -1188 3681 1188
rect 3635 -1200 3681 -1188
rect 3753 1188 3799 1200
rect 3753 -1188 3759 1188
rect 3793 -1188 3799 1188
rect 3753 -1200 3799 -1188
rect 3871 1188 3917 1200
rect 3871 -1188 3877 1188
rect 3911 -1188 3917 1188
rect 3871 -1200 3917 -1188
rect 3989 1188 4035 1200
rect 3989 -1188 3995 1188
rect 4029 -1188 4035 1188
rect 3989 -1200 4035 -1188
rect 4107 1188 4153 1200
rect 4107 -1188 4113 1188
rect 4147 -1188 4153 1188
rect 4107 -1200 4153 -1188
rect 4225 1188 4271 1200
rect 4225 -1188 4231 1188
rect 4265 -1188 4271 1188
rect 4225 -1200 4271 -1188
rect 4343 1188 4389 1200
rect 4343 -1188 4349 1188
rect 4383 -1188 4389 1188
rect 4343 -1200 4389 -1188
rect 4461 1188 4507 1200
rect 4461 -1188 4467 1188
rect 4501 -1188 4507 1188
rect 4461 -1200 4507 -1188
rect 4579 1188 4625 1200
rect 4579 -1188 4585 1188
rect 4619 -1188 4625 1188
rect 4579 -1200 4625 -1188
rect 4697 1188 4743 1200
rect 4697 -1188 4703 1188
rect 4737 -1188 4743 1188
rect 4697 -1200 4743 -1188
rect 4815 1188 4861 1200
rect 4815 -1188 4821 1188
rect 4855 -1188 4861 1188
rect 4815 -1200 4861 -1188
rect 4933 1188 4979 1200
rect 4933 -1188 4939 1188
rect 4973 -1188 4979 1188
rect 4933 -1200 4979 -1188
rect 5051 1188 5097 1200
rect 5051 -1188 5057 1188
rect 5091 -1188 5097 1188
rect 5051 -1200 5097 -1188
rect 5169 1188 5215 1200
rect 5169 -1188 5175 1188
rect 5209 -1188 5215 1188
rect 5169 -1200 5215 -1188
rect 5287 1188 5333 1200
rect 5287 -1188 5293 1188
rect 5327 -1188 5333 1188
rect 5287 -1200 5333 -1188
rect -5280 -1238 -5222 -1232
rect -5280 -1272 -5268 -1238
rect -5234 -1272 -5222 -1238
rect -5280 -1278 -5222 -1272
rect -5162 -1238 -5104 -1232
rect -5162 -1272 -5150 -1238
rect -5116 -1272 -5104 -1238
rect -5162 -1278 -5104 -1272
rect -5044 -1238 -4986 -1232
rect -5044 -1272 -5032 -1238
rect -4998 -1272 -4986 -1238
rect -5044 -1278 -4986 -1272
rect -4926 -1238 -4868 -1232
rect -4926 -1272 -4914 -1238
rect -4880 -1272 -4868 -1238
rect -4926 -1278 -4868 -1272
rect -4808 -1238 -4750 -1232
rect -4808 -1272 -4796 -1238
rect -4762 -1272 -4750 -1238
rect -4808 -1278 -4750 -1272
rect -4690 -1238 -4632 -1232
rect -4690 -1272 -4678 -1238
rect -4644 -1272 -4632 -1238
rect -4690 -1278 -4632 -1272
rect -4572 -1238 -4514 -1232
rect -4572 -1272 -4560 -1238
rect -4526 -1272 -4514 -1238
rect -4572 -1278 -4514 -1272
rect -4454 -1238 -4396 -1232
rect -4454 -1272 -4442 -1238
rect -4408 -1272 -4396 -1238
rect -4454 -1278 -4396 -1272
rect -4336 -1238 -4278 -1232
rect -4336 -1272 -4324 -1238
rect -4290 -1272 -4278 -1238
rect -4336 -1278 -4278 -1272
rect -4218 -1238 -4160 -1232
rect -4218 -1272 -4206 -1238
rect -4172 -1272 -4160 -1238
rect -4218 -1278 -4160 -1272
rect -4100 -1238 -4042 -1232
rect -4100 -1272 -4088 -1238
rect -4054 -1272 -4042 -1238
rect -4100 -1278 -4042 -1272
rect -3982 -1238 -3924 -1232
rect -3982 -1272 -3970 -1238
rect -3936 -1272 -3924 -1238
rect -3982 -1278 -3924 -1272
rect -3864 -1238 -3806 -1232
rect -3864 -1272 -3852 -1238
rect -3818 -1272 -3806 -1238
rect -3864 -1278 -3806 -1272
rect -3746 -1238 -3688 -1232
rect -3746 -1272 -3734 -1238
rect -3700 -1272 -3688 -1238
rect -3746 -1278 -3688 -1272
rect -3628 -1238 -3570 -1232
rect -3628 -1272 -3616 -1238
rect -3582 -1272 -3570 -1238
rect -3628 -1278 -3570 -1272
rect -3510 -1238 -3452 -1232
rect -3510 -1272 -3498 -1238
rect -3464 -1272 -3452 -1238
rect -3510 -1278 -3452 -1272
rect -3392 -1238 -3334 -1232
rect -3392 -1272 -3380 -1238
rect -3346 -1272 -3334 -1238
rect -3392 -1278 -3334 -1272
rect -3274 -1238 -3216 -1232
rect -3274 -1272 -3262 -1238
rect -3228 -1272 -3216 -1238
rect -3274 -1278 -3216 -1272
rect -3156 -1238 -3098 -1232
rect -3156 -1272 -3144 -1238
rect -3110 -1272 -3098 -1238
rect -3156 -1278 -3098 -1272
rect -3038 -1238 -2980 -1232
rect -3038 -1272 -3026 -1238
rect -2992 -1272 -2980 -1238
rect -3038 -1278 -2980 -1272
rect -2920 -1238 -2862 -1232
rect -2920 -1272 -2908 -1238
rect -2874 -1272 -2862 -1238
rect -2920 -1278 -2862 -1272
rect -2802 -1238 -2744 -1232
rect -2802 -1272 -2790 -1238
rect -2756 -1272 -2744 -1238
rect -2802 -1278 -2744 -1272
rect -2684 -1238 -2626 -1232
rect -2684 -1272 -2672 -1238
rect -2638 -1272 -2626 -1238
rect -2684 -1278 -2626 -1272
rect -2566 -1238 -2508 -1232
rect -2566 -1272 -2554 -1238
rect -2520 -1272 -2508 -1238
rect -2566 -1278 -2508 -1272
rect -2448 -1238 -2390 -1232
rect -2448 -1272 -2436 -1238
rect -2402 -1272 -2390 -1238
rect -2448 -1278 -2390 -1272
rect -2330 -1238 -2272 -1232
rect -2330 -1272 -2318 -1238
rect -2284 -1272 -2272 -1238
rect -2330 -1278 -2272 -1272
rect -2212 -1238 -2154 -1232
rect -2212 -1272 -2200 -1238
rect -2166 -1272 -2154 -1238
rect -2212 -1278 -2154 -1272
rect -2094 -1238 -2036 -1232
rect -2094 -1272 -2082 -1238
rect -2048 -1272 -2036 -1238
rect -2094 -1278 -2036 -1272
rect -1976 -1238 -1918 -1232
rect -1976 -1272 -1964 -1238
rect -1930 -1272 -1918 -1238
rect -1976 -1278 -1918 -1272
rect -1858 -1238 -1800 -1232
rect -1858 -1272 -1846 -1238
rect -1812 -1272 -1800 -1238
rect -1858 -1278 -1800 -1272
rect -1740 -1238 -1682 -1232
rect -1740 -1272 -1728 -1238
rect -1694 -1272 -1682 -1238
rect -1740 -1278 -1682 -1272
rect -1622 -1238 -1564 -1232
rect -1622 -1272 -1610 -1238
rect -1576 -1272 -1564 -1238
rect -1622 -1278 -1564 -1272
rect -1504 -1238 -1446 -1232
rect -1504 -1272 -1492 -1238
rect -1458 -1272 -1446 -1238
rect -1504 -1278 -1446 -1272
rect -1386 -1238 -1328 -1232
rect -1386 -1272 -1374 -1238
rect -1340 -1272 -1328 -1238
rect -1386 -1278 -1328 -1272
rect -1268 -1238 -1210 -1232
rect -1268 -1272 -1256 -1238
rect -1222 -1272 -1210 -1238
rect -1268 -1278 -1210 -1272
rect -1150 -1238 -1092 -1232
rect -1150 -1272 -1138 -1238
rect -1104 -1272 -1092 -1238
rect -1150 -1278 -1092 -1272
rect -1032 -1238 -974 -1232
rect -1032 -1272 -1020 -1238
rect -986 -1272 -974 -1238
rect -1032 -1278 -974 -1272
rect -914 -1238 -856 -1232
rect -914 -1272 -902 -1238
rect -868 -1272 -856 -1238
rect -914 -1278 -856 -1272
rect -796 -1238 -738 -1232
rect -796 -1272 -784 -1238
rect -750 -1272 -738 -1238
rect -796 -1278 -738 -1272
rect -678 -1238 -620 -1232
rect -678 -1272 -666 -1238
rect -632 -1272 -620 -1238
rect -678 -1278 -620 -1272
rect -560 -1238 -502 -1232
rect -560 -1272 -548 -1238
rect -514 -1272 -502 -1238
rect -560 -1278 -502 -1272
rect -442 -1238 -384 -1232
rect -442 -1272 -430 -1238
rect -396 -1272 -384 -1238
rect -442 -1278 -384 -1272
rect -324 -1238 -266 -1232
rect -324 -1272 -312 -1238
rect -278 -1272 -266 -1238
rect -324 -1278 -266 -1272
rect -206 -1238 -148 -1232
rect -206 -1272 -194 -1238
rect -160 -1272 -148 -1238
rect -206 -1278 -148 -1272
rect -88 -1238 -30 -1232
rect -88 -1272 -76 -1238
rect -42 -1272 -30 -1238
rect -88 -1278 -30 -1272
rect 30 -1238 88 -1232
rect 30 -1272 42 -1238
rect 76 -1272 88 -1238
rect 30 -1278 88 -1272
rect 148 -1238 206 -1232
rect 148 -1272 160 -1238
rect 194 -1272 206 -1238
rect 148 -1278 206 -1272
rect 266 -1238 324 -1232
rect 266 -1272 278 -1238
rect 312 -1272 324 -1238
rect 266 -1278 324 -1272
rect 384 -1238 442 -1232
rect 384 -1272 396 -1238
rect 430 -1272 442 -1238
rect 384 -1278 442 -1272
rect 502 -1238 560 -1232
rect 502 -1272 514 -1238
rect 548 -1272 560 -1238
rect 502 -1278 560 -1272
rect 620 -1238 678 -1232
rect 620 -1272 632 -1238
rect 666 -1272 678 -1238
rect 620 -1278 678 -1272
rect 738 -1238 796 -1232
rect 738 -1272 750 -1238
rect 784 -1272 796 -1238
rect 738 -1278 796 -1272
rect 856 -1238 914 -1232
rect 856 -1272 868 -1238
rect 902 -1272 914 -1238
rect 856 -1278 914 -1272
rect 974 -1238 1032 -1232
rect 974 -1272 986 -1238
rect 1020 -1272 1032 -1238
rect 974 -1278 1032 -1272
rect 1092 -1238 1150 -1232
rect 1092 -1272 1104 -1238
rect 1138 -1272 1150 -1238
rect 1092 -1278 1150 -1272
rect 1210 -1238 1268 -1232
rect 1210 -1272 1222 -1238
rect 1256 -1272 1268 -1238
rect 1210 -1278 1268 -1272
rect 1328 -1238 1386 -1232
rect 1328 -1272 1340 -1238
rect 1374 -1272 1386 -1238
rect 1328 -1278 1386 -1272
rect 1446 -1238 1504 -1232
rect 1446 -1272 1458 -1238
rect 1492 -1272 1504 -1238
rect 1446 -1278 1504 -1272
rect 1564 -1238 1622 -1232
rect 1564 -1272 1576 -1238
rect 1610 -1272 1622 -1238
rect 1564 -1278 1622 -1272
rect 1682 -1238 1740 -1232
rect 1682 -1272 1694 -1238
rect 1728 -1272 1740 -1238
rect 1682 -1278 1740 -1272
rect 1800 -1238 1858 -1232
rect 1800 -1272 1812 -1238
rect 1846 -1272 1858 -1238
rect 1800 -1278 1858 -1272
rect 1918 -1238 1976 -1232
rect 1918 -1272 1930 -1238
rect 1964 -1272 1976 -1238
rect 1918 -1278 1976 -1272
rect 2036 -1238 2094 -1232
rect 2036 -1272 2048 -1238
rect 2082 -1272 2094 -1238
rect 2036 -1278 2094 -1272
rect 2154 -1238 2212 -1232
rect 2154 -1272 2166 -1238
rect 2200 -1272 2212 -1238
rect 2154 -1278 2212 -1272
rect 2272 -1238 2330 -1232
rect 2272 -1272 2284 -1238
rect 2318 -1272 2330 -1238
rect 2272 -1278 2330 -1272
rect 2390 -1238 2448 -1232
rect 2390 -1272 2402 -1238
rect 2436 -1272 2448 -1238
rect 2390 -1278 2448 -1272
rect 2508 -1238 2566 -1232
rect 2508 -1272 2520 -1238
rect 2554 -1272 2566 -1238
rect 2508 -1278 2566 -1272
rect 2626 -1238 2684 -1232
rect 2626 -1272 2638 -1238
rect 2672 -1272 2684 -1238
rect 2626 -1278 2684 -1272
rect 2744 -1238 2802 -1232
rect 2744 -1272 2756 -1238
rect 2790 -1272 2802 -1238
rect 2744 -1278 2802 -1272
rect 2862 -1238 2920 -1232
rect 2862 -1272 2874 -1238
rect 2908 -1272 2920 -1238
rect 2862 -1278 2920 -1272
rect 2980 -1238 3038 -1232
rect 2980 -1272 2992 -1238
rect 3026 -1272 3038 -1238
rect 2980 -1278 3038 -1272
rect 3098 -1238 3156 -1232
rect 3098 -1272 3110 -1238
rect 3144 -1272 3156 -1238
rect 3098 -1278 3156 -1272
rect 3216 -1238 3274 -1232
rect 3216 -1272 3228 -1238
rect 3262 -1272 3274 -1238
rect 3216 -1278 3274 -1272
rect 3334 -1238 3392 -1232
rect 3334 -1272 3346 -1238
rect 3380 -1272 3392 -1238
rect 3334 -1278 3392 -1272
rect 3452 -1238 3510 -1232
rect 3452 -1272 3464 -1238
rect 3498 -1272 3510 -1238
rect 3452 -1278 3510 -1272
rect 3570 -1238 3628 -1232
rect 3570 -1272 3582 -1238
rect 3616 -1272 3628 -1238
rect 3570 -1278 3628 -1272
rect 3688 -1238 3746 -1232
rect 3688 -1272 3700 -1238
rect 3734 -1272 3746 -1238
rect 3688 -1278 3746 -1272
rect 3806 -1238 3864 -1232
rect 3806 -1272 3818 -1238
rect 3852 -1272 3864 -1238
rect 3806 -1278 3864 -1272
rect 3924 -1238 3982 -1232
rect 3924 -1272 3936 -1238
rect 3970 -1272 3982 -1238
rect 3924 -1278 3982 -1272
rect 4042 -1238 4100 -1232
rect 4042 -1272 4054 -1238
rect 4088 -1272 4100 -1238
rect 4042 -1278 4100 -1272
rect 4160 -1238 4218 -1232
rect 4160 -1272 4172 -1238
rect 4206 -1272 4218 -1238
rect 4160 -1278 4218 -1272
rect 4278 -1238 4336 -1232
rect 4278 -1272 4290 -1238
rect 4324 -1272 4336 -1238
rect 4278 -1278 4336 -1272
rect 4396 -1238 4454 -1232
rect 4396 -1272 4408 -1238
rect 4442 -1272 4454 -1238
rect 4396 -1278 4454 -1272
rect 4514 -1238 4572 -1232
rect 4514 -1272 4526 -1238
rect 4560 -1272 4572 -1238
rect 4514 -1278 4572 -1272
rect 4632 -1238 4690 -1232
rect 4632 -1272 4644 -1238
rect 4678 -1272 4690 -1238
rect 4632 -1278 4690 -1272
rect 4750 -1238 4808 -1232
rect 4750 -1272 4762 -1238
rect 4796 -1272 4808 -1238
rect 4750 -1278 4808 -1272
rect 4868 -1238 4926 -1232
rect 4868 -1272 4880 -1238
rect 4914 -1272 4926 -1238
rect 4868 -1278 4926 -1272
rect 4986 -1238 5044 -1232
rect 4986 -1272 4998 -1238
rect 5032 -1272 5044 -1238
rect 4986 -1278 5044 -1272
rect 5104 -1238 5162 -1232
rect 5104 -1272 5116 -1238
rect 5150 -1272 5162 -1238
rect 5104 -1278 5162 -1272
rect 5222 -1238 5280 -1232
rect 5222 -1272 5234 -1238
rect 5268 -1272 5280 -1238
rect 5222 -1278 5280 -1272
<< properties >>
string FIXED_BBOX -5424 -1357 5424 1357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 12 l 0.3 m 1 nf 90 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
