magic
tech sky130A
magscale 1 2
timestamp 1723380300
<< error_p >>
rect -3510 981 -3452 987
rect -3392 981 -3334 987
rect -3274 981 -3216 987
rect -3156 981 -3098 987
rect -3038 981 -2980 987
rect -2920 981 -2862 987
rect -2802 981 -2744 987
rect -2684 981 -2626 987
rect -2566 981 -2508 987
rect -2448 981 -2390 987
rect -2330 981 -2272 987
rect -2212 981 -2154 987
rect -2094 981 -2036 987
rect -1976 981 -1918 987
rect -1858 981 -1800 987
rect -1740 981 -1682 987
rect -1622 981 -1564 987
rect -1504 981 -1446 987
rect -1386 981 -1328 987
rect -1268 981 -1210 987
rect -1150 981 -1092 987
rect -1032 981 -974 987
rect -914 981 -856 987
rect -796 981 -738 987
rect -678 981 -620 987
rect -560 981 -502 987
rect -442 981 -384 987
rect -324 981 -266 987
rect -206 981 -148 987
rect -88 981 -30 987
rect 30 981 88 987
rect 148 981 206 987
rect 266 981 324 987
rect 384 981 442 987
rect 502 981 560 987
rect 620 981 678 987
rect 738 981 796 987
rect 856 981 914 987
rect 974 981 1032 987
rect 1092 981 1150 987
rect 1210 981 1268 987
rect 1328 981 1386 987
rect 1446 981 1504 987
rect 1564 981 1622 987
rect 1682 981 1740 987
rect 1800 981 1858 987
rect 1918 981 1976 987
rect 2036 981 2094 987
rect 2154 981 2212 987
rect 2272 981 2330 987
rect 2390 981 2448 987
rect 2508 981 2566 987
rect 2626 981 2684 987
rect 2744 981 2802 987
rect 2862 981 2920 987
rect 2980 981 3038 987
rect 3098 981 3156 987
rect 3216 981 3274 987
rect 3334 981 3392 987
rect 3452 981 3510 987
rect -3510 947 -3498 981
rect -3392 947 -3380 981
rect -3274 947 -3262 981
rect -3156 947 -3144 981
rect -3038 947 -3026 981
rect -2920 947 -2908 981
rect -2802 947 -2790 981
rect -2684 947 -2672 981
rect -2566 947 -2554 981
rect -2448 947 -2436 981
rect -2330 947 -2318 981
rect -2212 947 -2200 981
rect -2094 947 -2082 981
rect -1976 947 -1964 981
rect -1858 947 -1846 981
rect -1740 947 -1728 981
rect -1622 947 -1610 981
rect -1504 947 -1492 981
rect -1386 947 -1374 981
rect -1268 947 -1256 981
rect -1150 947 -1138 981
rect -1032 947 -1020 981
rect -914 947 -902 981
rect -796 947 -784 981
rect -678 947 -666 981
rect -560 947 -548 981
rect -442 947 -430 981
rect -324 947 -312 981
rect -206 947 -194 981
rect -88 947 -76 981
rect 30 947 42 981
rect 148 947 160 981
rect 266 947 278 981
rect 384 947 396 981
rect 502 947 514 981
rect 620 947 632 981
rect 738 947 750 981
rect 856 947 868 981
rect 974 947 986 981
rect 1092 947 1104 981
rect 1210 947 1222 981
rect 1328 947 1340 981
rect 1446 947 1458 981
rect 1564 947 1576 981
rect 1682 947 1694 981
rect 1800 947 1812 981
rect 1918 947 1930 981
rect 2036 947 2048 981
rect 2154 947 2166 981
rect 2272 947 2284 981
rect 2390 947 2402 981
rect 2508 947 2520 981
rect 2626 947 2638 981
rect 2744 947 2756 981
rect 2862 947 2874 981
rect 2980 947 2992 981
rect 3098 947 3110 981
rect 3216 947 3228 981
rect 3334 947 3346 981
rect 3452 947 3464 981
rect -3510 941 -3452 947
rect -3392 941 -3334 947
rect -3274 941 -3216 947
rect -3156 941 -3098 947
rect -3038 941 -2980 947
rect -2920 941 -2862 947
rect -2802 941 -2744 947
rect -2684 941 -2626 947
rect -2566 941 -2508 947
rect -2448 941 -2390 947
rect -2330 941 -2272 947
rect -2212 941 -2154 947
rect -2094 941 -2036 947
rect -1976 941 -1918 947
rect -1858 941 -1800 947
rect -1740 941 -1682 947
rect -1622 941 -1564 947
rect -1504 941 -1446 947
rect -1386 941 -1328 947
rect -1268 941 -1210 947
rect -1150 941 -1092 947
rect -1032 941 -974 947
rect -914 941 -856 947
rect -796 941 -738 947
rect -678 941 -620 947
rect -560 941 -502 947
rect -442 941 -384 947
rect -324 941 -266 947
rect -206 941 -148 947
rect -88 941 -30 947
rect 30 941 88 947
rect 148 941 206 947
rect 266 941 324 947
rect 384 941 442 947
rect 502 941 560 947
rect 620 941 678 947
rect 738 941 796 947
rect 856 941 914 947
rect 974 941 1032 947
rect 1092 941 1150 947
rect 1210 941 1268 947
rect 1328 941 1386 947
rect 1446 941 1504 947
rect 1564 941 1622 947
rect 1682 941 1740 947
rect 1800 941 1858 947
rect 1918 941 1976 947
rect 2036 941 2094 947
rect 2154 941 2212 947
rect 2272 941 2330 947
rect 2390 941 2448 947
rect 2508 941 2566 947
rect 2626 941 2684 947
rect 2744 941 2802 947
rect 2862 941 2920 947
rect 2980 941 3038 947
rect 3098 941 3156 947
rect 3216 941 3274 947
rect 3334 941 3392 947
rect 3452 941 3510 947
rect -3510 -947 -3452 -941
rect -3392 -947 -3334 -941
rect -3274 -947 -3216 -941
rect -3156 -947 -3098 -941
rect -3038 -947 -2980 -941
rect -2920 -947 -2862 -941
rect -2802 -947 -2744 -941
rect -2684 -947 -2626 -941
rect -2566 -947 -2508 -941
rect -2448 -947 -2390 -941
rect -2330 -947 -2272 -941
rect -2212 -947 -2154 -941
rect -2094 -947 -2036 -941
rect -1976 -947 -1918 -941
rect -1858 -947 -1800 -941
rect -1740 -947 -1682 -941
rect -1622 -947 -1564 -941
rect -1504 -947 -1446 -941
rect -1386 -947 -1328 -941
rect -1268 -947 -1210 -941
rect -1150 -947 -1092 -941
rect -1032 -947 -974 -941
rect -914 -947 -856 -941
rect -796 -947 -738 -941
rect -678 -947 -620 -941
rect -560 -947 -502 -941
rect -442 -947 -384 -941
rect -324 -947 -266 -941
rect -206 -947 -148 -941
rect -88 -947 -30 -941
rect 30 -947 88 -941
rect 148 -947 206 -941
rect 266 -947 324 -941
rect 384 -947 442 -941
rect 502 -947 560 -941
rect 620 -947 678 -941
rect 738 -947 796 -941
rect 856 -947 914 -941
rect 974 -947 1032 -941
rect 1092 -947 1150 -941
rect 1210 -947 1268 -941
rect 1328 -947 1386 -941
rect 1446 -947 1504 -941
rect 1564 -947 1622 -941
rect 1682 -947 1740 -941
rect 1800 -947 1858 -941
rect 1918 -947 1976 -941
rect 2036 -947 2094 -941
rect 2154 -947 2212 -941
rect 2272 -947 2330 -941
rect 2390 -947 2448 -941
rect 2508 -947 2566 -941
rect 2626 -947 2684 -941
rect 2744 -947 2802 -941
rect 2862 -947 2920 -941
rect 2980 -947 3038 -941
rect 3098 -947 3156 -941
rect 3216 -947 3274 -941
rect 3334 -947 3392 -941
rect 3452 -947 3510 -941
rect -3510 -981 -3498 -947
rect -3392 -981 -3380 -947
rect -3274 -981 -3262 -947
rect -3156 -981 -3144 -947
rect -3038 -981 -3026 -947
rect -2920 -981 -2908 -947
rect -2802 -981 -2790 -947
rect -2684 -981 -2672 -947
rect -2566 -981 -2554 -947
rect -2448 -981 -2436 -947
rect -2330 -981 -2318 -947
rect -2212 -981 -2200 -947
rect -2094 -981 -2082 -947
rect -1976 -981 -1964 -947
rect -1858 -981 -1846 -947
rect -1740 -981 -1728 -947
rect -1622 -981 -1610 -947
rect -1504 -981 -1492 -947
rect -1386 -981 -1374 -947
rect -1268 -981 -1256 -947
rect -1150 -981 -1138 -947
rect -1032 -981 -1020 -947
rect -914 -981 -902 -947
rect -796 -981 -784 -947
rect -678 -981 -666 -947
rect -560 -981 -548 -947
rect -442 -981 -430 -947
rect -324 -981 -312 -947
rect -206 -981 -194 -947
rect -88 -981 -76 -947
rect 30 -981 42 -947
rect 148 -981 160 -947
rect 266 -981 278 -947
rect 384 -981 396 -947
rect 502 -981 514 -947
rect 620 -981 632 -947
rect 738 -981 750 -947
rect 856 -981 868 -947
rect 974 -981 986 -947
rect 1092 -981 1104 -947
rect 1210 -981 1222 -947
rect 1328 -981 1340 -947
rect 1446 -981 1458 -947
rect 1564 -981 1576 -947
rect 1682 -981 1694 -947
rect 1800 -981 1812 -947
rect 1918 -981 1930 -947
rect 2036 -981 2048 -947
rect 2154 -981 2166 -947
rect 2272 -981 2284 -947
rect 2390 -981 2402 -947
rect 2508 -981 2520 -947
rect 2626 -981 2638 -947
rect 2744 -981 2756 -947
rect 2862 -981 2874 -947
rect 2980 -981 2992 -947
rect 3098 -981 3110 -947
rect 3216 -981 3228 -947
rect 3334 -981 3346 -947
rect 3452 -981 3464 -947
rect -3510 -987 -3452 -981
rect -3392 -987 -3334 -981
rect -3274 -987 -3216 -981
rect -3156 -987 -3098 -981
rect -3038 -987 -2980 -981
rect -2920 -987 -2862 -981
rect -2802 -987 -2744 -981
rect -2684 -987 -2626 -981
rect -2566 -987 -2508 -981
rect -2448 -987 -2390 -981
rect -2330 -987 -2272 -981
rect -2212 -987 -2154 -981
rect -2094 -987 -2036 -981
rect -1976 -987 -1918 -981
rect -1858 -987 -1800 -981
rect -1740 -987 -1682 -981
rect -1622 -987 -1564 -981
rect -1504 -987 -1446 -981
rect -1386 -987 -1328 -981
rect -1268 -987 -1210 -981
rect -1150 -987 -1092 -981
rect -1032 -987 -974 -981
rect -914 -987 -856 -981
rect -796 -987 -738 -981
rect -678 -987 -620 -981
rect -560 -987 -502 -981
rect -442 -987 -384 -981
rect -324 -987 -266 -981
rect -206 -987 -148 -981
rect -88 -987 -30 -981
rect 30 -987 88 -981
rect 148 -987 206 -981
rect 266 -987 324 -981
rect 384 -987 442 -981
rect 502 -987 560 -981
rect 620 -987 678 -981
rect 738 -987 796 -981
rect 856 -987 914 -981
rect 974 -987 1032 -981
rect 1092 -987 1150 -981
rect 1210 -987 1268 -981
rect 1328 -987 1386 -981
rect 1446 -987 1504 -981
rect 1564 -987 1622 -981
rect 1682 -987 1740 -981
rect 1800 -987 1858 -981
rect 1918 -987 1976 -981
rect 2036 -987 2094 -981
rect 2154 -987 2212 -981
rect 2272 -987 2330 -981
rect 2390 -987 2448 -981
rect 2508 -987 2566 -981
rect 2626 -987 2684 -981
rect 2744 -987 2802 -981
rect 2862 -987 2920 -981
rect 2980 -987 3038 -981
rect 3098 -987 3156 -981
rect 3216 -987 3274 -981
rect 3334 -987 3392 -981
rect 3452 -987 3510 -981
<< nwell >>
rect -3707 -1119 3707 1119
<< pmos >>
rect -3511 -900 -3451 900
rect -3393 -900 -3333 900
rect -3275 -900 -3215 900
rect -3157 -900 -3097 900
rect -3039 -900 -2979 900
rect -2921 -900 -2861 900
rect -2803 -900 -2743 900
rect -2685 -900 -2625 900
rect -2567 -900 -2507 900
rect -2449 -900 -2389 900
rect -2331 -900 -2271 900
rect -2213 -900 -2153 900
rect -2095 -900 -2035 900
rect -1977 -900 -1917 900
rect -1859 -900 -1799 900
rect -1741 -900 -1681 900
rect -1623 -900 -1563 900
rect -1505 -900 -1445 900
rect -1387 -900 -1327 900
rect -1269 -900 -1209 900
rect -1151 -900 -1091 900
rect -1033 -900 -973 900
rect -915 -900 -855 900
rect -797 -900 -737 900
rect -679 -900 -619 900
rect -561 -900 -501 900
rect -443 -900 -383 900
rect -325 -900 -265 900
rect -207 -900 -147 900
rect -89 -900 -29 900
rect 29 -900 89 900
rect 147 -900 207 900
rect 265 -900 325 900
rect 383 -900 443 900
rect 501 -900 561 900
rect 619 -900 679 900
rect 737 -900 797 900
rect 855 -900 915 900
rect 973 -900 1033 900
rect 1091 -900 1151 900
rect 1209 -900 1269 900
rect 1327 -900 1387 900
rect 1445 -900 1505 900
rect 1563 -900 1623 900
rect 1681 -900 1741 900
rect 1799 -900 1859 900
rect 1917 -900 1977 900
rect 2035 -900 2095 900
rect 2153 -900 2213 900
rect 2271 -900 2331 900
rect 2389 -900 2449 900
rect 2507 -900 2567 900
rect 2625 -900 2685 900
rect 2743 -900 2803 900
rect 2861 -900 2921 900
rect 2979 -900 3039 900
rect 3097 -900 3157 900
rect 3215 -900 3275 900
rect 3333 -900 3393 900
rect 3451 -900 3511 900
<< pdiff >>
rect -3569 888 -3511 900
rect -3569 -888 -3557 888
rect -3523 -888 -3511 888
rect -3569 -900 -3511 -888
rect -3451 888 -3393 900
rect -3451 -888 -3439 888
rect -3405 -888 -3393 888
rect -3451 -900 -3393 -888
rect -3333 888 -3275 900
rect -3333 -888 -3321 888
rect -3287 -888 -3275 888
rect -3333 -900 -3275 -888
rect -3215 888 -3157 900
rect -3215 -888 -3203 888
rect -3169 -888 -3157 888
rect -3215 -900 -3157 -888
rect -3097 888 -3039 900
rect -3097 -888 -3085 888
rect -3051 -888 -3039 888
rect -3097 -900 -3039 -888
rect -2979 888 -2921 900
rect -2979 -888 -2967 888
rect -2933 -888 -2921 888
rect -2979 -900 -2921 -888
rect -2861 888 -2803 900
rect -2861 -888 -2849 888
rect -2815 -888 -2803 888
rect -2861 -900 -2803 -888
rect -2743 888 -2685 900
rect -2743 -888 -2731 888
rect -2697 -888 -2685 888
rect -2743 -900 -2685 -888
rect -2625 888 -2567 900
rect -2625 -888 -2613 888
rect -2579 -888 -2567 888
rect -2625 -900 -2567 -888
rect -2507 888 -2449 900
rect -2507 -888 -2495 888
rect -2461 -888 -2449 888
rect -2507 -900 -2449 -888
rect -2389 888 -2331 900
rect -2389 -888 -2377 888
rect -2343 -888 -2331 888
rect -2389 -900 -2331 -888
rect -2271 888 -2213 900
rect -2271 -888 -2259 888
rect -2225 -888 -2213 888
rect -2271 -900 -2213 -888
rect -2153 888 -2095 900
rect -2153 -888 -2141 888
rect -2107 -888 -2095 888
rect -2153 -900 -2095 -888
rect -2035 888 -1977 900
rect -2035 -888 -2023 888
rect -1989 -888 -1977 888
rect -2035 -900 -1977 -888
rect -1917 888 -1859 900
rect -1917 -888 -1905 888
rect -1871 -888 -1859 888
rect -1917 -900 -1859 -888
rect -1799 888 -1741 900
rect -1799 -888 -1787 888
rect -1753 -888 -1741 888
rect -1799 -900 -1741 -888
rect -1681 888 -1623 900
rect -1681 -888 -1669 888
rect -1635 -888 -1623 888
rect -1681 -900 -1623 -888
rect -1563 888 -1505 900
rect -1563 -888 -1551 888
rect -1517 -888 -1505 888
rect -1563 -900 -1505 -888
rect -1445 888 -1387 900
rect -1445 -888 -1433 888
rect -1399 -888 -1387 888
rect -1445 -900 -1387 -888
rect -1327 888 -1269 900
rect -1327 -888 -1315 888
rect -1281 -888 -1269 888
rect -1327 -900 -1269 -888
rect -1209 888 -1151 900
rect -1209 -888 -1197 888
rect -1163 -888 -1151 888
rect -1209 -900 -1151 -888
rect -1091 888 -1033 900
rect -1091 -888 -1079 888
rect -1045 -888 -1033 888
rect -1091 -900 -1033 -888
rect -973 888 -915 900
rect -973 -888 -961 888
rect -927 -888 -915 888
rect -973 -900 -915 -888
rect -855 888 -797 900
rect -855 -888 -843 888
rect -809 -888 -797 888
rect -855 -900 -797 -888
rect -737 888 -679 900
rect -737 -888 -725 888
rect -691 -888 -679 888
rect -737 -900 -679 -888
rect -619 888 -561 900
rect -619 -888 -607 888
rect -573 -888 -561 888
rect -619 -900 -561 -888
rect -501 888 -443 900
rect -501 -888 -489 888
rect -455 -888 -443 888
rect -501 -900 -443 -888
rect -383 888 -325 900
rect -383 -888 -371 888
rect -337 -888 -325 888
rect -383 -900 -325 -888
rect -265 888 -207 900
rect -265 -888 -253 888
rect -219 -888 -207 888
rect -265 -900 -207 -888
rect -147 888 -89 900
rect -147 -888 -135 888
rect -101 -888 -89 888
rect -147 -900 -89 -888
rect -29 888 29 900
rect -29 -888 -17 888
rect 17 -888 29 888
rect -29 -900 29 -888
rect 89 888 147 900
rect 89 -888 101 888
rect 135 -888 147 888
rect 89 -900 147 -888
rect 207 888 265 900
rect 207 -888 219 888
rect 253 -888 265 888
rect 207 -900 265 -888
rect 325 888 383 900
rect 325 -888 337 888
rect 371 -888 383 888
rect 325 -900 383 -888
rect 443 888 501 900
rect 443 -888 455 888
rect 489 -888 501 888
rect 443 -900 501 -888
rect 561 888 619 900
rect 561 -888 573 888
rect 607 -888 619 888
rect 561 -900 619 -888
rect 679 888 737 900
rect 679 -888 691 888
rect 725 -888 737 888
rect 679 -900 737 -888
rect 797 888 855 900
rect 797 -888 809 888
rect 843 -888 855 888
rect 797 -900 855 -888
rect 915 888 973 900
rect 915 -888 927 888
rect 961 -888 973 888
rect 915 -900 973 -888
rect 1033 888 1091 900
rect 1033 -888 1045 888
rect 1079 -888 1091 888
rect 1033 -900 1091 -888
rect 1151 888 1209 900
rect 1151 -888 1163 888
rect 1197 -888 1209 888
rect 1151 -900 1209 -888
rect 1269 888 1327 900
rect 1269 -888 1281 888
rect 1315 -888 1327 888
rect 1269 -900 1327 -888
rect 1387 888 1445 900
rect 1387 -888 1399 888
rect 1433 -888 1445 888
rect 1387 -900 1445 -888
rect 1505 888 1563 900
rect 1505 -888 1517 888
rect 1551 -888 1563 888
rect 1505 -900 1563 -888
rect 1623 888 1681 900
rect 1623 -888 1635 888
rect 1669 -888 1681 888
rect 1623 -900 1681 -888
rect 1741 888 1799 900
rect 1741 -888 1753 888
rect 1787 -888 1799 888
rect 1741 -900 1799 -888
rect 1859 888 1917 900
rect 1859 -888 1871 888
rect 1905 -888 1917 888
rect 1859 -900 1917 -888
rect 1977 888 2035 900
rect 1977 -888 1989 888
rect 2023 -888 2035 888
rect 1977 -900 2035 -888
rect 2095 888 2153 900
rect 2095 -888 2107 888
rect 2141 -888 2153 888
rect 2095 -900 2153 -888
rect 2213 888 2271 900
rect 2213 -888 2225 888
rect 2259 -888 2271 888
rect 2213 -900 2271 -888
rect 2331 888 2389 900
rect 2331 -888 2343 888
rect 2377 -888 2389 888
rect 2331 -900 2389 -888
rect 2449 888 2507 900
rect 2449 -888 2461 888
rect 2495 -888 2507 888
rect 2449 -900 2507 -888
rect 2567 888 2625 900
rect 2567 -888 2579 888
rect 2613 -888 2625 888
rect 2567 -900 2625 -888
rect 2685 888 2743 900
rect 2685 -888 2697 888
rect 2731 -888 2743 888
rect 2685 -900 2743 -888
rect 2803 888 2861 900
rect 2803 -888 2815 888
rect 2849 -888 2861 888
rect 2803 -900 2861 -888
rect 2921 888 2979 900
rect 2921 -888 2933 888
rect 2967 -888 2979 888
rect 2921 -900 2979 -888
rect 3039 888 3097 900
rect 3039 -888 3051 888
rect 3085 -888 3097 888
rect 3039 -900 3097 -888
rect 3157 888 3215 900
rect 3157 -888 3169 888
rect 3203 -888 3215 888
rect 3157 -900 3215 -888
rect 3275 888 3333 900
rect 3275 -888 3287 888
rect 3321 -888 3333 888
rect 3275 -900 3333 -888
rect 3393 888 3451 900
rect 3393 -888 3405 888
rect 3439 -888 3451 888
rect 3393 -900 3451 -888
rect 3511 888 3569 900
rect 3511 -888 3523 888
rect 3557 -888 3569 888
rect 3511 -900 3569 -888
<< pdiffc >>
rect -3557 -888 -3523 888
rect -3439 -888 -3405 888
rect -3321 -888 -3287 888
rect -3203 -888 -3169 888
rect -3085 -888 -3051 888
rect -2967 -888 -2933 888
rect -2849 -888 -2815 888
rect -2731 -888 -2697 888
rect -2613 -888 -2579 888
rect -2495 -888 -2461 888
rect -2377 -888 -2343 888
rect -2259 -888 -2225 888
rect -2141 -888 -2107 888
rect -2023 -888 -1989 888
rect -1905 -888 -1871 888
rect -1787 -888 -1753 888
rect -1669 -888 -1635 888
rect -1551 -888 -1517 888
rect -1433 -888 -1399 888
rect -1315 -888 -1281 888
rect -1197 -888 -1163 888
rect -1079 -888 -1045 888
rect -961 -888 -927 888
rect -843 -888 -809 888
rect -725 -888 -691 888
rect -607 -888 -573 888
rect -489 -888 -455 888
rect -371 -888 -337 888
rect -253 -888 -219 888
rect -135 -888 -101 888
rect -17 -888 17 888
rect 101 -888 135 888
rect 219 -888 253 888
rect 337 -888 371 888
rect 455 -888 489 888
rect 573 -888 607 888
rect 691 -888 725 888
rect 809 -888 843 888
rect 927 -888 961 888
rect 1045 -888 1079 888
rect 1163 -888 1197 888
rect 1281 -888 1315 888
rect 1399 -888 1433 888
rect 1517 -888 1551 888
rect 1635 -888 1669 888
rect 1753 -888 1787 888
rect 1871 -888 1905 888
rect 1989 -888 2023 888
rect 2107 -888 2141 888
rect 2225 -888 2259 888
rect 2343 -888 2377 888
rect 2461 -888 2495 888
rect 2579 -888 2613 888
rect 2697 -888 2731 888
rect 2815 -888 2849 888
rect 2933 -888 2967 888
rect 3051 -888 3085 888
rect 3169 -888 3203 888
rect 3287 -888 3321 888
rect 3405 -888 3439 888
rect 3523 -888 3557 888
<< nsubdiff >>
rect -3671 1049 -3575 1083
rect 3575 1049 3671 1083
rect -3671 987 -3637 1049
rect 3637 987 3671 1049
rect -3671 -1049 -3637 -987
rect 3637 -1049 3671 -987
rect -3671 -1083 -3575 -1049
rect 3575 -1083 3671 -1049
<< nsubdiffcont >>
rect -3575 1049 3575 1083
rect -3671 -987 -3637 987
rect 3637 -987 3671 987
rect -3575 -1083 3575 -1049
<< poly >>
rect -3514 981 -3448 997
rect -3514 947 -3498 981
rect -3464 947 -3448 981
rect -3514 931 -3448 947
rect -3396 981 -3330 997
rect -3396 947 -3380 981
rect -3346 947 -3330 981
rect -3396 931 -3330 947
rect -3278 981 -3212 997
rect -3278 947 -3262 981
rect -3228 947 -3212 981
rect -3278 931 -3212 947
rect -3160 981 -3094 997
rect -3160 947 -3144 981
rect -3110 947 -3094 981
rect -3160 931 -3094 947
rect -3042 981 -2976 997
rect -3042 947 -3026 981
rect -2992 947 -2976 981
rect -3042 931 -2976 947
rect -2924 981 -2858 997
rect -2924 947 -2908 981
rect -2874 947 -2858 981
rect -2924 931 -2858 947
rect -2806 981 -2740 997
rect -2806 947 -2790 981
rect -2756 947 -2740 981
rect -2806 931 -2740 947
rect -2688 981 -2622 997
rect -2688 947 -2672 981
rect -2638 947 -2622 981
rect -2688 931 -2622 947
rect -2570 981 -2504 997
rect -2570 947 -2554 981
rect -2520 947 -2504 981
rect -2570 931 -2504 947
rect -2452 981 -2386 997
rect -2452 947 -2436 981
rect -2402 947 -2386 981
rect -2452 931 -2386 947
rect -2334 981 -2268 997
rect -2334 947 -2318 981
rect -2284 947 -2268 981
rect -2334 931 -2268 947
rect -2216 981 -2150 997
rect -2216 947 -2200 981
rect -2166 947 -2150 981
rect -2216 931 -2150 947
rect -2098 981 -2032 997
rect -2098 947 -2082 981
rect -2048 947 -2032 981
rect -2098 931 -2032 947
rect -1980 981 -1914 997
rect -1980 947 -1964 981
rect -1930 947 -1914 981
rect -1980 931 -1914 947
rect -1862 981 -1796 997
rect -1862 947 -1846 981
rect -1812 947 -1796 981
rect -1862 931 -1796 947
rect -1744 981 -1678 997
rect -1744 947 -1728 981
rect -1694 947 -1678 981
rect -1744 931 -1678 947
rect -1626 981 -1560 997
rect -1626 947 -1610 981
rect -1576 947 -1560 981
rect -1626 931 -1560 947
rect -1508 981 -1442 997
rect -1508 947 -1492 981
rect -1458 947 -1442 981
rect -1508 931 -1442 947
rect -1390 981 -1324 997
rect -1390 947 -1374 981
rect -1340 947 -1324 981
rect -1390 931 -1324 947
rect -1272 981 -1206 997
rect -1272 947 -1256 981
rect -1222 947 -1206 981
rect -1272 931 -1206 947
rect -1154 981 -1088 997
rect -1154 947 -1138 981
rect -1104 947 -1088 981
rect -1154 931 -1088 947
rect -1036 981 -970 997
rect -1036 947 -1020 981
rect -986 947 -970 981
rect -1036 931 -970 947
rect -918 981 -852 997
rect -918 947 -902 981
rect -868 947 -852 981
rect -918 931 -852 947
rect -800 981 -734 997
rect -800 947 -784 981
rect -750 947 -734 981
rect -800 931 -734 947
rect -682 981 -616 997
rect -682 947 -666 981
rect -632 947 -616 981
rect -682 931 -616 947
rect -564 981 -498 997
rect -564 947 -548 981
rect -514 947 -498 981
rect -564 931 -498 947
rect -446 981 -380 997
rect -446 947 -430 981
rect -396 947 -380 981
rect -446 931 -380 947
rect -328 981 -262 997
rect -328 947 -312 981
rect -278 947 -262 981
rect -328 931 -262 947
rect -210 981 -144 997
rect -210 947 -194 981
rect -160 947 -144 981
rect -210 931 -144 947
rect -92 981 -26 997
rect -92 947 -76 981
rect -42 947 -26 981
rect -92 931 -26 947
rect 26 981 92 997
rect 26 947 42 981
rect 76 947 92 981
rect 26 931 92 947
rect 144 981 210 997
rect 144 947 160 981
rect 194 947 210 981
rect 144 931 210 947
rect 262 981 328 997
rect 262 947 278 981
rect 312 947 328 981
rect 262 931 328 947
rect 380 981 446 997
rect 380 947 396 981
rect 430 947 446 981
rect 380 931 446 947
rect 498 981 564 997
rect 498 947 514 981
rect 548 947 564 981
rect 498 931 564 947
rect 616 981 682 997
rect 616 947 632 981
rect 666 947 682 981
rect 616 931 682 947
rect 734 981 800 997
rect 734 947 750 981
rect 784 947 800 981
rect 734 931 800 947
rect 852 981 918 997
rect 852 947 868 981
rect 902 947 918 981
rect 852 931 918 947
rect 970 981 1036 997
rect 970 947 986 981
rect 1020 947 1036 981
rect 970 931 1036 947
rect 1088 981 1154 997
rect 1088 947 1104 981
rect 1138 947 1154 981
rect 1088 931 1154 947
rect 1206 981 1272 997
rect 1206 947 1222 981
rect 1256 947 1272 981
rect 1206 931 1272 947
rect 1324 981 1390 997
rect 1324 947 1340 981
rect 1374 947 1390 981
rect 1324 931 1390 947
rect 1442 981 1508 997
rect 1442 947 1458 981
rect 1492 947 1508 981
rect 1442 931 1508 947
rect 1560 981 1626 997
rect 1560 947 1576 981
rect 1610 947 1626 981
rect 1560 931 1626 947
rect 1678 981 1744 997
rect 1678 947 1694 981
rect 1728 947 1744 981
rect 1678 931 1744 947
rect 1796 981 1862 997
rect 1796 947 1812 981
rect 1846 947 1862 981
rect 1796 931 1862 947
rect 1914 981 1980 997
rect 1914 947 1930 981
rect 1964 947 1980 981
rect 1914 931 1980 947
rect 2032 981 2098 997
rect 2032 947 2048 981
rect 2082 947 2098 981
rect 2032 931 2098 947
rect 2150 981 2216 997
rect 2150 947 2166 981
rect 2200 947 2216 981
rect 2150 931 2216 947
rect 2268 981 2334 997
rect 2268 947 2284 981
rect 2318 947 2334 981
rect 2268 931 2334 947
rect 2386 981 2452 997
rect 2386 947 2402 981
rect 2436 947 2452 981
rect 2386 931 2452 947
rect 2504 981 2570 997
rect 2504 947 2520 981
rect 2554 947 2570 981
rect 2504 931 2570 947
rect 2622 981 2688 997
rect 2622 947 2638 981
rect 2672 947 2688 981
rect 2622 931 2688 947
rect 2740 981 2806 997
rect 2740 947 2756 981
rect 2790 947 2806 981
rect 2740 931 2806 947
rect 2858 981 2924 997
rect 2858 947 2874 981
rect 2908 947 2924 981
rect 2858 931 2924 947
rect 2976 981 3042 997
rect 2976 947 2992 981
rect 3026 947 3042 981
rect 2976 931 3042 947
rect 3094 981 3160 997
rect 3094 947 3110 981
rect 3144 947 3160 981
rect 3094 931 3160 947
rect 3212 981 3278 997
rect 3212 947 3228 981
rect 3262 947 3278 981
rect 3212 931 3278 947
rect 3330 981 3396 997
rect 3330 947 3346 981
rect 3380 947 3396 981
rect 3330 931 3396 947
rect 3448 981 3514 997
rect 3448 947 3464 981
rect 3498 947 3514 981
rect 3448 931 3514 947
rect -3511 900 -3451 931
rect -3393 900 -3333 931
rect -3275 900 -3215 931
rect -3157 900 -3097 931
rect -3039 900 -2979 931
rect -2921 900 -2861 931
rect -2803 900 -2743 931
rect -2685 900 -2625 931
rect -2567 900 -2507 931
rect -2449 900 -2389 931
rect -2331 900 -2271 931
rect -2213 900 -2153 931
rect -2095 900 -2035 931
rect -1977 900 -1917 931
rect -1859 900 -1799 931
rect -1741 900 -1681 931
rect -1623 900 -1563 931
rect -1505 900 -1445 931
rect -1387 900 -1327 931
rect -1269 900 -1209 931
rect -1151 900 -1091 931
rect -1033 900 -973 931
rect -915 900 -855 931
rect -797 900 -737 931
rect -679 900 -619 931
rect -561 900 -501 931
rect -443 900 -383 931
rect -325 900 -265 931
rect -207 900 -147 931
rect -89 900 -29 931
rect 29 900 89 931
rect 147 900 207 931
rect 265 900 325 931
rect 383 900 443 931
rect 501 900 561 931
rect 619 900 679 931
rect 737 900 797 931
rect 855 900 915 931
rect 973 900 1033 931
rect 1091 900 1151 931
rect 1209 900 1269 931
rect 1327 900 1387 931
rect 1445 900 1505 931
rect 1563 900 1623 931
rect 1681 900 1741 931
rect 1799 900 1859 931
rect 1917 900 1977 931
rect 2035 900 2095 931
rect 2153 900 2213 931
rect 2271 900 2331 931
rect 2389 900 2449 931
rect 2507 900 2567 931
rect 2625 900 2685 931
rect 2743 900 2803 931
rect 2861 900 2921 931
rect 2979 900 3039 931
rect 3097 900 3157 931
rect 3215 900 3275 931
rect 3333 900 3393 931
rect 3451 900 3511 931
rect -3511 -931 -3451 -900
rect -3393 -931 -3333 -900
rect -3275 -931 -3215 -900
rect -3157 -931 -3097 -900
rect -3039 -931 -2979 -900
rect -2921 -931 -2861 -900
rect -2803 -931 -2743 -900
rect -2685 -931 -2625 -900
rect -2567 -931 -2507 -900
rect -2449 -931 -2389 -900
rect -2331 -931 -2271 -900
rect -2213 -931 -2153 -900
rect -2095 -931 -2035 -900
rect -1977 -931 -1917 -900
rect -1859 -931 -1799 -900
rect -1741 -931 -1681 -900
rect -1623 -931 -1563 -900
rect -1505 -931 -1445 -900
rect -1387 -931 -1327 -900
rect -1269 -931 -1209 -900
rect -1151 -931 -1091 -900
rect -1033 -931 -973 -900
rect -915 -931 -855 -900
rect -797 -931 -737 -900
rect -679 -931 -619 -900
rect -561 -931 -501 -900
rect -443 -931 -383 -900
rect -325 -931 -265 -900
rect -207 -931 -147 -900
rect -89 -931 -29 -900
rect 29 -931 89 -900
rect 147 -931 207 -900
rect 265 -931 325 -900
rect 383 -931 443 -900
rect 501 -931 561 -900
rect 619 -931 679 -900
rect 737 -931 797 -900
rect 855 -931 915 -900
rect 973 -931 1033 -900
rect 1091 -931 1151 -900
rect 1209 -931 1269 -900
rect 1327 -931 1387 -900
rect 1445 -931 1505 -900
rect 1563 -931 1623 -900
rect 1681 -931 1741 -900
rect 1799 -931 1859 -900
rect 1917 -931 1977 -900
rect 2035 -931 2095 -900
rect 2153 -931 2213 -900
rect 2271 -931 2331 -900
rect 2389 -931 2449 -900
rect 2507 -931 2567 -900
rect 2625 -931 2685 -900
rect 2743 -931 2803 -900
rect 2861 -931 2921 -900
rect 2979 -931 3039 -900
rect 3097 -931 3157 -900
rect 3215 -931 3275 -900
rect 3333 -931 3393 -900
rect 3451 -931 3511 -900
rect -3514 -947 -3448 -931
rect -3514 -981 -3498 -947
rect -3464 -981 -3448 -947
rect -3514 -997 -3448 -981
rect -3396 -947 -3330 -931
rect -3396 -981 -3380 -947
rect -3346 -981 -3330 -947
rect -3396 -997 -3330 -981
rect -3278 -947 -3212 -931
rect -3278 -981 -3262 -947
rect -3228 -981 -3212 -947
rect -3278 -997 -3212 -981
rect -3160 -947 -3094 -931
rect -3160 -981 -3144 -947
rect -3110 -981 -3094 -947
rect -3160 -997 -3094 -981
rect -3042 -947 -2976 -931
rect -3042 -981 -3026 -947
rect -2992 -981 -2976 -947
rect -3042 -997 -2976 -981
rect -2924 -947 -2858 -931
rect -2924 -981 -2908 -947
rect -2874 -981 -2858 -947
rect -2924 -997 -2858 -981
rect -2806 -947 -2740 -931
rect -2806 -981 -2790 -947
rect -2756 -981 -2740 -947
rect -2806 -997 -2740 -981
rect -2688 -947 -2622 -931
rect -2688 -981 -2672 -947
rect -2638 -981 -2622 -947
rect -2688 -997 -2622 -981
rect -2570 -947 -2504 -931
rect -2570 -981 -2554 -947
rect -2520 -981 -2504 -947
rect -2570 -997 -2504 -981
rect -2452 -947 -2386 -931
rect -2452 -981 -2436 -947
rect -2402 -981 -2386 -947
rect -2452 -997 -2386 -981
rect -2334 -947 -2268 -931
rect -2334 -981 -2318 -947
rect -2284 -981 -2268 -947
rect -2334 -997 -2268 -981
rect -2216 -947 -2150 -931
rect -2216 -981 -2200 -947
rect -2166 -981 -2150 -947
rect -2216 -997 -2150 -981
rect -2098 -947 -2032 -931
rect -2098 -981 -2082 -947
rect -2048 -981 -2032 -947
rect -2098 -997 -2032 -981
rect -1980 -947 -1914 -931
rect -1980 -981 -1964 -947
rect -1930 -981 -1914 -947
rect -1980 -997 -1914 -981
rect -1862 -947 -1796 -931
rect -1862 -981 -1846 -947
rect -1812 -981 -1796 -947
rect -1862 -997 -1796 -981
rect -1744 -947 -1678 -931
rect -1744 -981 -1728 -947
rect -1694 -981 -1678 -947
rect -1744 -997 -1678 -981
rect -1626 -947 -1560 -931
rect -1626 -981 -1610 -947
rect -1576 -981 -1560 -947
rect -1626 -997 -1560 -981
rect -1508 -947 -1442 -931
rect -1508 -981 -1492 -947
rect -1458 -981 -1442 -947
rect -1508 -997 -1442 -981
rect -1390 -947 -1324 -931
rect -1390 -981 -1374 -947
rect -1340 -981 -1324 -947
rect -1390 -997 -1324 -981
rect -1272 -947 -1206 -931
rect -1272 -981 -1256 -947
rect -1222 -981 -1206 -947
rect -1272 -997 -1206 -981
rect -1154 -947 -1088 -931
rect -1154 -981 -1138 -947
rect -1104 -981 -1088 -947
rect -1154 -997 -1088 -981
rect -1036 -947 -970 -931
rect -1036 -981 -1020 -947
rect -986 -981 -970 -947
rect -1036 -997 -970 -981
rect -918 -947 -852 -931
rect -918 -981 -902 -947
rect -868 -981 -852 -947
rect -918 -997 -852 -981
rect -800 -947 -734 -931
rect -800 -981 -784 -947
rect -750 -981 -734 -947
rect -800 -997 -734 -981
rect -682 -947 -616 -931
rect -682 -981 -666 -947
rect -632 -981 -616 -947
rect -682 -997 -616 -981
rect -564 -947 -498 -931
rect -564 -981 -548 -947
rect -514 -981 -498 -947
rect -564 -997 -498 -981
rect -446 -947 -380 -931
rect -446 -981 -430 -947
rect -396 -981 -380 -947
rect -446 -997 -380 -981
rect -328 -947 -262 -931
rect -328 -981 -312 -947
rect -278 -981 -262 -947
rect -328 -997 -262 -981
rect -210 -947 -144 -931
rect -210 -981 -194 -947
rect -160 -981 -144 -947
rect -210 -997 -144 -981
rect -92 -947 -26 -931
rect -92 -981 -76 -947
rect -42 -981 -26 -947
rect -92 -997 -26 -981
rect 26 -947 92 -931
rect 26 -981 42 -947
rect 76 -981 92 -947
rect 26 -997 92 -981
rect 144 -947 210 -931
rect 144 -981 160 -947
rect 194 -981 210 -947
rect 144 -997 210 -981
rect 262 -947 328 -931
rect 262 -981 278 -947
rect 312 -981 328 -947
rect 262 -997 328 -981
rect 380 -947 446 -931
rect 380 -981 396 -947
rect 430 -981 446 -947
rect 380 -997 446 -981
rect 498 -947 564 -931
rect 498 -981 514 -947
rect 548 -981 564 -947
rect 498 -997 564 -981
rect 616 -947 682 -931
rect 616 -981 632 -947
rect 666 -981 682 -947
rect 616 -997 682 -981
rect 734 -947 800 -931
rect 734 -981 750 -947
rect 784 -981 800 -947
rect 734 -997 800 -981
rect 852 -947 918 -931
rect 852 -981 868 -947
rect 902 -981 918 -947
rect 852 -997 918 -981
rect 970 -947 1036 -931
rect 970 -981 986 -947
rect 1020 -981 1036 -947
rect 970 -997 1036 -981
rect 1088 -947 1154 -931
rect 1088 -981 1104 -947
rect 1138 -981 1154 -947
rect 1088 -997 1154 -981
rect 1206 -947 1272 -931
rect 1206 -981 1222 -947
rect 1256 -981 1272 -947
rect 1206 -997 1272 -981
rect 1324 -947 1390 -931
rect 1324 -981 1340 -947
rect 1374 -981 1390 -947
rect 1324 -997 1390 -981
rect 1442 -947 1508 -931
rect 1442 -981 1458 -947
rect 1492 -981 1508 -947
rect 1442 -997 1508 -981
rect 1560 -947 1626 -931
rect 1560 -981 1576 -947
rect 1610 -981 1626 -947
rect 1560 -997 1626 -981
rect 1678 -947 1744 -931
rect 1678 -981 1694 -947
rect 1728 -981 1744 -947
rect 1678 -997 1744 -981
rect 1796 -947 1862 -931
rect 1796 -981 1812 -947
rect 1846 -981 1862 -947
rect 1796 -997 1862 -981
rect 1914 -947 1980 -931
rect 1914 -981 1930 -947
rect 1964 -981 1980 -947
rect 1914 -997 1980 -981
rect 2032 -947 2098 -931
rect 2032 -981 2048 -947
rect 2082 -981 2098 -947
rect 2032 -997 2098 -981
rect 2150 -947 2216 -931
rect 2150 -981 2166 -947
rect 2200 -981 2216 -947
rect 2150 -997 2216 -981
rect 2268 -947 2334 -931
rect 2268 -981 2284 -947
rect 2318 -981 2334 -947
rect 2268 -997 2334 -981
rect 2386 -947 2452 -931
rect 2386 -981 2402 -947
rect 2436 -981 2452 -947
rect 2386 -997 2452 -981
rect 2504 -947 2570 -931
rect 2504 -981 2520 -947
rect 2554 -981 2570 -947
rect 2504 -997 2570 -981
rect 2622 -947 2688 -931
rect 2622 -981 2638 -947
rect 2672 -981 2688 -947
rect 2622 -997 2688 -981
rect 2740 -947 2806 -931
rect 2740 -981 2756 -947
rect 2790 -981 2806 -947
rect 2740 -997 2806 -981
rect 2858 -947 2924 -931
rect 2858 -981 2874 -947
rect 2908 -981 2924 -947
rect 2858 -997 2924 -981
rect 2976 -947 3042 -931
rect 2976 -981 2992 -947
rect 3026 -981 3042 -947
rect 2976 -997 3042 -981
rect 3094 -947 3160 -931
rect 3094 -981 3110 -947
rect 3144 -981 3160 -947
rect 3094 -997 3160 -981
rect 3212 -947 3278 -931
rect 3212 -981 3228 -947
rect 3262 -981 3278 -947
rect 3212 -997 3278 -981
rect 3330 -947 3396 -931
rect 3330 -981 3346 -947
rect 3380 -981 3396 -947
rect 3330 -997 3396 -981
rect 3448 -947 3514 -931
rect 3448 -981 3464 -947
rect 3498 -981 3514 -947
rect 3448 -997 3514 -981
<< polycont >>
rect -3498 947 -3464 981
rect -3380 947 -3346 981
rect -3262 947 -3228 981
rect -3144 947 -3110 981
rect -3026 947 -2992 981
rect -2908 947 -2874 981
rect -2790 947 -2756 981
rect -2672 947 -2638 981
rect -2554 947 -2520 981
rect -2436 947 -2402 981
rect -2318 947 -2284 981
rect -2200 947 -2166 981
rect -2082 947 -2048 981
rect -1964 947 -1930 981
rect -1846 947 -1812 981
rect -1728 947 -1694 981
rect -1610 947 -1576 981
rect -1492 947 -1458 981
rect -1374 947 -1340 981
rect -1256 947 -1222 981
rect -1138 947 -1104 981
rect -1020 947 -986 981
rect -902 947 -868 981
rect -784 947 -750 981
rect -666 947 -632 981
rect -548 947 -514 981
rect -430 947 -396 981
rect -312 947 -278 981
rect -194 947 -160 981
rect -76 947 -42 981
rect 42 947 76 981
rect 160 947 194 981
rect 278 947 312 981
rect 396 947 430 981
rect 514 947 548 981
rect 632 947 666 981
rect 750 947 784 981
rect 868 947 902 981
rect 986 947 1020 981
rect 1104 947 1138 981
rect 1222 947 1256 981
rect 1340 947 1374 981
rect 1458 947 1492 981
rect 1576 947 1610 981
rect 1694 947 1728 981
rect 1812 947 1846 981
rect 1930 947 1964 981
rect 2048 947 2082 981
rect 2166 947 2200 981
rect 2284 947 2318 981
rect 2402 947 2436 981
rect 2520 947 2554 981
rect 2638 947 2672 981
rect 2756 947 2790 981
rect 2874 947 2908 981
rect 2992 947 3026 981
rect 3110 947 3144 981
rect 3228 947 3262 981
rect 3346 947 3380 981
rect 3464 947 3498 981
rect -3498 -981 -3464 -947
rect -3380 -981 -3346 -947
rect -3262 -981 -3228 -947
rect -3144 -981 -3110 -947
rect -3026 -981 -2992 -947
rect -2908 -981 -2874 -947
rect -2790 -981 -2756 -947
rect -2672 -981 -2638 -947
rect -2554 -981 -2520 -947
rect -2436 -981 -2402 -947
rect -2318 -981 -2284 -947
rect -2200 -981 -2166 -947
rect -2082 -981 -2048 -947
rect -1964 -981 -1930 -947
rect -1846 -981 -1812 -947
rect -1728 -981 -1694 -947
rect -1610 -981 -1576 -947
rect -1492 -981 -1458 -947
rect -1374 -981 -1340 -947
rect -1256 -981 -1222 -947
rect -1138 -981 -1104 -947
rect -1020 -981 -986 -947
rect -902 -981 -868 -947
rect -784 -981 -750 -947
rect -666 -981 -632 -947
rect -548 -981 -514 -947
rect -430 -981 -396 -947
rect -312 -981 -278 -947
rect -194 -981 -160 -947
rect -76 -981 -42 -947
rect 42 -981 76 -947
rect 160 -981 194 -947
rect 278 -981 312 -947
rect 396 -981 430 -947
rect 514 -981 548 -947
rect 632 -981 666 -947
rect 750 -981 784 -947
rect 868 -981 902 -947
rect 986 -981 1020 -947
rect 1104 -981 1138 -947
rect 1222 -981 1256 -947
rect 1340 -981 1374 -947
rect 1458 -981 1492 -947
rect 1576 -981 1610 -947
rect 1694 -981 1728 -947
rect 1812 -981 1846 -947
rect 1930 -981 1964 -947
rect 2048 -981 2082 -947
rect 2166 -981 2200 -947
rect 2284 -981 2318 -947
rect 2402 -981 2436 -947
rect 2520 -981 2554 -947
rect 2638 -981 2672 -947
rect 2756 -981 2790 -947
rect 2874 -981 2908 -947
rect 2992 -981 3026 -947
rect 3110 -981 3144 -947
rect 3228 -981 3262 -947
rect 3346 -981 3380 -947
rect 3464 -981 3498 -947
<< locali >>
rect -3671 1049 -3575 1083
rect 3575 1049 3671 1083
rect -3671 987 -3637 1049
rect 3637 987 3671 1049
rect -3514 947 -3498 981
rect -3464 947 -3448 981
rect -3396 947 -3380 981
rect -3346 947 -3330 981
rect -3278 947 -3262 981
rect -3228 947 -3212 981
rect -3160 947 -3144 981
rect -3110 947 -3094 981
rect -3042 947 -3026 981
rect -2992 947 -2976 981
rect -2924 947 -2908 981
rect -2874 947 -2858 981
rect -2806 947 -2790 981
rect -2756 947 -2740 981
rect -2688 947 -2672 981
rect -2638 947 -2622 981
rect -2570 947 -2554 981
rect -2520 947 -2504 981
rect -2452 947 -2436 981
rect -2402 947 -2386 981
rect -2334 947 -2318 981
rect -2284 947 -2268 981
rect -2216 947 -2200 981
rect -2166 947 -2150 981
rect -2098 947 -2082 981
rect -2048 947 -2032 981
rect -1980 947 -1964 981
rect -1930 947 -1914 981
rect -1862 947 -1846 981
rect -1812 947 -1796 981
rect -1744 947 -1728 981
rect -1694 947 -1678 981
rect -1626 947 -1610 981
rect -1576 947 -1560 981
rect -1508 947 -1492 981
rect -1458 947 -1442 981
rect -1390 947 -1374 981
rect -1340 947 -1324 981
rect -1272 947 -1256 981
rect -1222 947 -1206 981
rect -1154 947 -1138 981
rect -1104 947 -1088 981
rect -1036 947 -1020 981
rect -986 947 -970 981
rect -918 947 -902 981
rect -868 947 -852 981
rect -800 947 -784 981
rect -750 947 -734 981
rect -682 947 -666 981
rect -632 947 -616 981
rect -564 947 -548 981
rect -514 947 -498 981
rect -446 947 -430 981
rect -396 947 -380 981
rect -328 947 -312 981
rect -278 947 -262 981
rect -210 947 -194 981
rect -160 947 -144 981
rect -92 947 -76 981
rect -42 947 -26 981
rect 26 947 42 981
rect 76 947 92 981
rect 144 947 160 981
rect 194 947 210 981
rect 262 947 278 981
rect 312 947 328 981
rect 380 947 396 981
rect 430 947 446 981
rect 498 947 514 981
rect 548 947 564 981
rect 616 947 632 981
rect 666 947 682 981
rect 734 947 750 981
rect 784 947 800 981
rect 852 947 868 981
rect 902 947 918 981
rect 970 947 986 981
rect 1020 947 1036 981
rect 1088 947 1104 981
rect 1138 947 1154 981
rect 1206 947 1222 981
rect 1256 947 1272 981
rect 1324 947 1340 981
rect 1374 947 1390 981
rect 1442 947 1458 981
rect 1492 947 1508 981
rect 1560 947 1576 981
rect 1610 947 1626 981
rect 1678 947 1694 981
rect 1728 947 1744 981
rect 1796 947 1812 981
rect 1846 947 1862 981
rect 1914 947 1930 981
rect 1964 947 1980 981
rect 2032 947 2048 981
rect 2082 947 2098 981
rect 2150 947 2166 981
rect 2200 947 2216 981
rect 2268 947 2284 981
rect 2318 947 2334 981
rect 2386 947 2402 981
rect 2436 947 2452 981
rect 2504 947 2520 981
rect 2554 947 2570 981
rect 2622 947 2638 981
rect 2672 947 2688 981
rect 2740 947 2756 981
rect 2790 947 2806 981
rect 2858 947 2874 981
rect 2908 947 2924 981
rect 2976 947 2992 981
rect 3026 947 3042 981
rect 3094 947 3110 981
rect 3144 947 3160 981
rect 3212 947 3228 981
rect 3262 947 3278 981
rect 3330 947 3346 981
rect 3380 947 3396 981
rect 3448 947 3464 981
rect 3498 947 3514 981
rect -3557 888 -3523 904
rect -3557 -904 -3523 -888
rect -3439 888 -3405 904
rect -3439 -904 -3405 -888
rect -3321 888 -3287 904
rect -3321 -904 -3287 -888
rect -3203 888 -3169 904
rect -3203 -904 -3169 -888
rect -3085 888 -3051 904
rect -3085 -904 -3051 -888
rect -2967 888 -2933 904
rect -2967 -904 -2933 -888
rect -2849 888 -2815 904
rect -2849 -904 -2815 -888
rect -2731 888 -2697 904
rect -2731 -904 -2697 -888
rect -2613 888 -2579 904
rect -2613 -904 -2579 -888
rect -2495 888 -2461 904
rect -2495 -904 -2461 -888
rect -2377 888 -2343 904
rect -2377 -904 -2343 -888
rect -2259 888 -2225 904
rect -2259 -904 -2225 -888
rect -2141 888 -2107 904
rect -2141 -904 -2107 -888
rect -2023 888 -1989 904
rect -2023 -904 -1989 -888
rect -1905 888 -1871 904
rect -1905 -904 -1871 -888
rect -1787 888 -1753 904
rect -1787 -904 -1753 -888
rect -1669 888 -1635 904
rect -1669 -904 -1635 -888
rect -1551 888 -1517 904
rect -1551 -904 -1517 -888
rect -1433 888 -1399 904
rect -1433 -904 -1399 -888
rect -1315 888 -1281 904
rect -1315 -904 -1281 -888
rect -1197 888 -1163 904
rect -1197 -904 -1163 -888
rect -1079 888 -1045 904
rect -1079 -904 -1045 -888
rect -961 888 -927 904
rect -961 -904 -927 -888
rect -843 888 -809 904
rect -843 -904 -809 -888
rect -725 888 -691 904
rect -725 -904 -691 -888
rect -607 888 -573 904
rect -607 -904 -573 -888
rect -489 888 -455 904
rect -489 -904 -455 -888
rect -371 888 -337 904
rect -371 -904 -337 -888
rect -253 888 -219 904
rect -253 -904 -219 -888
rect -135 888 -101 904
rect -135 -904 -101 -888
rect -17 888 17 904
rect -17 -904 17 -888
rect 101 888 135 904
rect 101 -904 135 -888
rect 219 888 253 904
rect 219 -904 253 -888
rect 337 888 371 904
rect 337 -904 371 -888
rect 455 888 489 904
rect 455 -904 489 -888
rect 573 888 607 904
rect 573 -904 607 -888
rect 691 888 725 904
rect 691 -904 725 -888
rect 809 888 843 904
rect 809 -904 843 -888
rect 927 888 961 904
rect 927 -904 961 -888
rect 1045 888 1079 904
rect 1045 -904 1079 -888
rect 1163 888 1197 904
rect 1163 -904 1197 -888
rect 1281 888 1315 904
rect 1281 -904 1315 -888
rect 1399 888 1433 904
rect 1399 -904 1433 -888
rect 1517 888 1551 904
rect 1517 -904 1551 -888
rect 1635 888 1669 904
rect 1635 -904 1669 -888
rect 1753 888 1787 904
rect 1753 -904 1787 -888
rect 1871 888 1905 904
rect 1871 -904 1905 -888
rect 1989 888 2023 904
rect 1989 -904 2023 -888
rect 2107 888 2141 904
rect 2107 -904 2141 -888
rect 2225 888 2259 904
rect 2225 -904 2259 -888
rect 2343 888 2377 904
rect 2343 -904 2377 -888
rect 2461 888 2495 904
rect 2461 -904 2495 -888
rect 2579 888 2613 904
rect 2579 -904 2613 -888
rect 2697 888 2731 904
rect 2697 -904 2731 -888
rect 2815 888 2849 904
rect 2815 -904 2849 -888
rect 2933 888 2967 904
rect 2933 -904 2967 -888
rect 3051 888 3085 904
rect 3051 -904 3085 -888
rect 3169 888 3203 904
rect 3169 -904 3203 -888
rect 3287 888 3321 904
rect 3287 -904 3321 -888
rect 3405 888 3439 904
rect 3405 -904 3439 -888
rect 3523 888 3557 904
rect 3523 -904 3557 -888
rect -3514 -981 -3498 -947
rect -3464 -981 -3448 -947
rect -3396 -981 -3380 -947
rect -3346 -981 -3330 -947
rect -3278 -981 -3262 -947
rect -3228 -981 -3212 -947
rect -3160 -981 -3144 -947
rect -3110 -981 -3094 -947
rect -3042 -981 -3026 -947
rect -2992 -981 -2976 -947
rect -2924 -981 -2908 -947
rect -2874 -981 -2858 -947
rect -2806 -981 -2790 -947
rect -2756 -981 -2740 -947
rect -2688 -981 -2672 -947
rect -2638 -981 -2622 -947
rect -2570 -981 -2554 -947
rect -2520 -981 -2504 -947
rect -2452 -981 -2436 -947
rect -2402 -981 -2386 -947
rect -2334 -981 -2318 -947
rect -2284 -981 -2268 -947
rect -2216 -981 -2200 -947
rect -2166 -981 -2150 -947
rect -2098 -981 -2082 -947
rect -2048 -981 -2032 -947
rect -1980 -981 -1964 -947
rect -1930 -981 -1914 -947
rect -1862 -981 -1846 -947
rect -1812 -981 -1796 -947
rect -1744 -981 -1728 -947
rect -1694 -981 -1678 -947
rect -1626 -981 -1610 -947
rect -1576 -981 -1560 -947
rect -1508 -981 -1492 -947
rect -1458 -981 -1442 -947
rect -1390 -981 -1374 -947
rect -1340 -981 -1324 -947
rect -1272 -981 -1256 -947
rect -1222 -981 -1206 -947
rect -1154 -981 -1138 -947
rect -1104 -981 -1088 -947
rect -1036 -981 -1020 -947
rect -986 -981 -970 -947
rect -918 -981 -902 -947
rect -868 -981 -852 -947
rect -800 -981 -784 -947
rect -750 -981 -734 -947
rect -682 -981 -666 -947
rect -632 -981 -616 -947
rect -564 -981 -548 -947
rect -514 -981 -498 -947
rect -446 -981 -430 -947
rect -396 -981 -380 -947
rect -328 -981 -312 -947
rect -278 -981 -262 -947
rect -210 -981 -194 -947
rect -160 -981 -144 -947
rect -92 -981 -76 -947
rect -42 -981 -26 -947
rect 26 -981 42 -947
rect 76 -981 92 -947
rect 144 -981 160 -947
rect 194 -981 210 -947
rect 262 -981 278 -947
rect 312 -981 328 -947
rect 380 -981 396 -947
rect 430 -981 446 -947
rect 498 -981 514 -947
rect 548 -981 564 -947
rect 616 -981 632 -947
rect 666 -981 682 -947
rect 734 -981 750 -947
rect 784 -981 800 -947
rect 852 -981 868 -947
rect 902 -981 918 -947
rect 970 -981 986 -947
rect 1020 -981 1036 -947
rect 1088 -981 1104 -947
rect 1138 -981 1154 -947
rect 1206 -981 1222 -947
rect 1256 -981 1272 -947
rect 1324 -981 1340 -947
rect 1374 -981 1390 -947
rect 1442 -981 1458 -947
rect 1492 -981 1508 -947
rect 1560 -981 1576 -947
rect 1610 -981 1626 -947
rect 1678 -981 1694 -947
rect 1728 -981 1744 -947
rect 1796 -981 1812 -947
rect 1846 -981 1862 -947
rect 1914 -981 1930 -947
rect 1964 -981 1980 -947
rect 2032 -981 2048 -947
rect 2082 -981 2098 -947
rect 2150 -981 2166 -947
rect 2200 -981 2216 -947
rect 2268 -981 2284 -947
rect 2318 -981 2334 -947
rect 2386 -981 2402 -947
rect 2436 -981 2452 -947
rect 2504 -981 2520 -947
rect 2554 -981 2570 -947
rect 2622 -981 2638 -947
rect 2672 -981 2688 -947
rect 2740 -981 2756 -947
rect 2790 -981 2806 -947
rect 2858 -981 2874 -947
rect 2908 -981 2924 -947
rect 2976 -981 2992 -947
rect 3026 -981 3042 -947
rect 3094 -981 3110 -947
rect 3144 -981 3160 -947
rect 3212 -981 3228 -947
rect 3262 -981 3278 -947
rect 3330 -981 3346 -947
rect 3380 -981 3396 -947
rect 3448 -981 3464 -947
rect 3498 -981 3514 -947
rect -3671 -1049 -3637 -987
rect 3637 -1049 3671 -987
rect -3671 -1083 -3575 -1049
rect 3575 -1083 3671 -1049
<< viali >>
rect -3498 947 -3464 981
rect -3380 947 -3346 981
rect -3262 947 -3228 981
rect -3144 947 -3110 981
rect -3026 947 -2992 981
rect -2908 947 -2874 981
rect -2790 947 -2756 981
rect -2672 947 -2638 981
rect -2554 947 -2520 981
rect -2436 947 -2402 981
rect -2318 947 -2284 981
rect -2200 947 -2166 981
rect -2082 947 -2048 981
rect -1964 947 -1930 981
rect -1846 947 -1812 981
rect -1728 947 -1694 981
rect -1610 947 -1576 981
rect -1492 947 -1458 981
rect -1374 947 -1340 981
rect -1256 947 -1222 981
rect -1138 947 -1104 981
rect -1020 947 -986 981
rect -902 947 -868 981
rect -784 947 -750 981
rect -666 947 -632 981
rect -548 947 -514 981
rect -430 947 -396 981
rect -312 947 -278 981
rect -194 947 -160 981
rect -76 947 -42 981
rect 42 947 76 981
rect 160 947 194 981
rect 278 947 312 981
rect 396 947 430 981
rect 514 947 548 981
rect 632 947 666 981
rect 750 947 784 981
rect 868 947 902 981
rect 986 947 1020 981
rect 1104 947 1138 981
rect 1222 947 1256 981
rect 1340 947 1374 981
rect 1458 947 1492 981
rect 1576 947 1610 981
rect 1694 947 1728 981
rect 1812 947 1846 981
rect 1930 947 1964 981
rect 2048 947 2082 981
rect 2166 947 2200 981
rect 2284 947 2318 981
rect 2402 947 2436 981
rect 2520 947 2554 981
rect 2638 947 2672 981
rect 2756 947 2790 981
rect 2874 947 2908 981
rect 2992 947 3026 981
rect 3110 947 3144 981
rect 3228 947 3262 981
rect 3346 947 3380 981
rect 3464 947 3498 981
rect -3557 -888 -3523 888
rect -3439 -888 -3405 888
rect -3321 -888 -3287 888
rect -3203 -888 -3169 888
rect -3085 -888 -3051 888
rect -2967 -888 -2933 888
rect -2849 -888 -2815 888
rect -2731 -888 -2697 888
rect -2613 -888 -2579 888
rect -2495 -888 -2461 888
rect -2377 -888 -2343 888
rect -2259 -888 -2225 888
rect -2141 -888 -2107 888
rect -2023 -888 -1989 888
rect -1905 -888 -1871 888
rect -1787 -888 -1753 888
rect -1669 -888 -1635 888
rect -1551 -888 -1517 888
rect -1433 -888 -1399 888
rect -1315 -888 -1281 888
rect -1197 -888 -1163 888
rect -1079 -888 -1045 888
rect -961 -888 -927 888
rect -843 -888 -809 888
rect -725 -888 -691 888
rect -607 -888 -573 888
rect -489 -888 -455 888
rect -371 -888 -337 888
rect -253 -888 -219 888
rect -135 -888 -101 888
rect -17 -888 17 888
rect 101 -888 135 888
rect 219 -888 253 888
rect 337 -888 371 888
rect 455 -888 489 888
rect 573 -888 607 888
rect 691 -888 725 888
rect 809 -888 843 888
rect 927 -888 961 888
rect 1045 -888 1079 888
rect 1163 -888 1197 888
rect 1281 -888 1315 888
rect 1399 -888 1433 888
rect 1517 -888 1551 888
rect 1635 -888 1669 888
rect 1753 -888 1787 888
rect 1871 -888 1905 888
rect 1989 -888 2023 888
rect 2107 -888 2141 888
rect 2225 -888 2259 888
rect 2343 -888 2377 888
rect 2461 -888 2495 888
rect 2579 -888 2613 888
rect 2697 -888 2731 888
rect 2815 -888 2849 888
rect 2933 -888 2967 888
rect 3051 -888 3085 888
rect 3169 -888 3203 888
rect 3287 -888 3321 888
rect 3405 -888 3439 888
rect 3523 -888 3557 888
rect -3498 -981 -3464 -947
rect -3380 -981 -3346 -947
rect -3262 -981 -3228 -947
rect -3144 -981 -3110 -947
rect -3026 -981 -2992 -947
rect -2908 -981 -2874 -947
rect -2790 -981 -2756 -947
rect -2672 -981 -2638 -947
rect -2554 -981 -2520 -947
rect -2436 -981 -2402 -947
rect -2318 -981 -2284 -947
rect -2200 -981 -2166 -947
rect -2082 -981 -2048 -947
rect -1964 -981 -1930 -947
rect -1846 -981 -1812 -947
rect -1728 -981 -1694 -947
rect -1610 -981 -1576 -947
rect -1492 -981 -1458 -947
rect -1374 -981 -1340 -947
rect -1256 -981 -1222 -947
rect -1138 -981 -1104 -947
rect -1020 -981 -986 -947
rect -902 -981 -868 -947
rect -784 -981 -750 -947
rect -666 -981 -632 -947
rect -548 -981 -514 -947
rect -430 -981 -396 -947
rect -312 -981 -278 -947
rect -194 -981 -160 -947
rect -76 -981 -42 -947
rect 42 -981 76 -947
rect 160 -981 194 -947
rect 278 -981 312 -947
rect 396 -981 430 -947
rect 514 -981 548 -947
rect 632 -981 666 -947
rect 750 -981 784 -947
rect 868 -981 902 -947
rect 986 -981 1020 -947
rect 1104 -981 1138 -947
rect 1222 -981 1256 -947
rect 1340 -981 1374 -947
rect 1458 -981 1492 -947
rect 1576 -981 1610 -947
rect 1694 -981 1728 -947
rect 1812 -981 1846 -947
rect 1930 -981 1964 -947
rect 2048 -981 2082 -947
rect 2166 -981 2200 -947
rect 2284 -981 2318 -947
rect 2402 -981 2436 -947
rect 2520 -981 2554 -947
rect 2638 -981 2672 -947
rect 2756 -981 2790 -947
rect 2874 -981 2908 -947
rect 2992 -981 3026 -947
rect 3110 -981 3144 -947
rect 3228 -981 3262 -947
rect 3346 -981 3380 -947
rect 3464 -981 3498 -947
<< metal1 >>
rect -3510 981 -3452 987
rect -3510 947 -3498 981
rect -3464 947 -3452 981
rect -3510 941 -3452 947
rect -3392 981 -3334 987
rect -3392 947 -3380 981
rect -3346 947 -3334 981
rect -3392 941 -3334 947
rect -3274 981 -3216 987
rect -3274 947 -3262 981
rect -3228 947 -3216 981
rect -3274 941 -3216 947
rect -3156 981 -3098 987
rect -3156 947 -3144 981
rect -3110 947 -3098 981
rect -3156 941 -3098 947
rect -3038 981 -2980 987
rect -3038 947 -3026 981
rect -2992 947 -2980 981
rect -3038 941 -2980 947
rect -2920 981 -2862 987
rect -2920 947 -2908 981
rect -2874 947 -2862 981
rect -2920 941 -2862 947
rect -2802 981 -2744 987
rect -2802 947 -2790 981
rect -2756 947 -2744 981
rect -2802 941 -2744 947
rect -2684 981 -2626 987
rect -2684 947 -2672 981
rect -2638 947 -2626 981
rect -2684 941 -2626 947
rect -2566 981 -2508 987
rect -2566 947 -2554 981
rect -2520 947 -2508 981
rect -2566 941 -2508 947
rect -2448 981 -2390 987
rect -2448 947 -2436 981
rect -2402 947 -2390 981
rect -2448 941 -2390 947
rect -2330 981 -2272 987
rect -2330 947 -2318 981
rect -2284 947 -2272 981
rect -2330 941 -2272 947
rect -2212 981 -2154 987
rect -2212 947 -2200 981
rect -2166 947 -2154 981
rect -2212 941 -2154 947
rect -2094 981 -2036 987
rect -2094 947 -2082 981
rect -2048 947 -2036 981
rect -2094 941 -2036 947
rect -1976 981 -1918 987
rect -1976 947 -1964 981
rect -1930 947 -1918 981
rect -1976 941 -1918 947
rect -1858 981 -1800 987
rect -1858 947 -1846 981
rect -1812 947 -1800 981
rect -1858 941 -1800 947
rect -1740 981 -1682 987
rect -1740 947 -1728 981
rect -1694 947 -1682 981
rect -1740 941 -1682 947
rect -1622 981 -1564 987
rect -1622 947 -1610 981
rect -1576 947 -1564 981
rect -1622 941 -1564 947
rect -1504 981 -1446 987
rect -1504 947 -1492 981
rect -1458 947 -1446 981
rect -1504 941 -1446 947
rect -1386 981 -1328 987
rect -1386 947 -1374 981
rect -1340 947 -1328 981
rect -1386 941 -1328 947
rect -1268 981 -1210 987
rect -1268 947 -1256 981
rect -1222 947 -1210 981
rect -1268 941 -1210 947
rect -1150 981 -1092 987
rect -1150 947 -1138 981
rect -1104 947 -1092 981
rect -1150 941 -1092 947
rect -1032 981 -974 987
rect -1032 947 -1020 981
rect -986 947 -974 981
rect -1032 941 -974 947
rect -914 981 -856 987
rect -914 947 -902 981
rect -868 947 -856 981
rect -914 941 -856 947
rect -796 981 -738 987
rect -796 947 -784 981
rect -750 947 -738 981
rect -796 941 -738 947
rect -678 981 -620 987
rect -678 947 -666 981
rect -632 947 -620 981
rect -678 941 -620 947
rect -560 981 -502 987
rect -560 947 -548 981
rect -514 947 -502 981
rect -560 941 -502 947
rect -442 981 -384 987
rect -442 947 -430 981
rect -396 947 -384 981
rect -442 941 -384 947
rect -324 981 -266 987
rect -324 947 -312 981
rect -278 947 -266 981
rect -324 941 -266 947
rect -206 981 -148 987
rect -206 947 -194 981
rect -160 947 -148 981
rect -206 941 -148 947
rect -88 981 -30 987
rect -88 947 -76 981
rect -42 947 -30 981
rect -88 941 -30 947
rect 30 981 88 987
rect 30 947 42 981
rect 76 947 88 981
rect 30 941 88 947
rect 148 981 206 987
rect 148 947 160 981
rect 194 947 206 981
rect 148 941 206 947
rect 266 981 324 987
rect 266 947 278 981
rect 312 947 324 981
rect 266 941 324 947
rect 384 981 442 987
rect 384 947 396 981
rect 430 947 442 981
rect 384 941 442 947
rect 502 981 560 987
rect 502 947 514 981
rect 548 947 560 981
rect 502 941 560 947
rect 620 981 678 987
rect 620 947 632 981
rect 666 947 678 981
rect 620 941 678 947
rect 738 981 796 987
rect 738 947 750 981
rect 784 947 796 981
rect 738 941 796 947
rect 856 981 914 987
rect 856 947 868 981
rect 902 947 914 981
rect 856 941 914 947
rect 974 981 1032 987
rect 974 947 986 981
rect 1020 947 1032 981
rect 974 941 1032 947
rect 1092 981 1150 987
rect 1092 947 1104 981
rect 1138 947 1150 981
rect 1092 941 1150 947
rect 1210 981 1268 987
rect 1210 947 1222 981
rect 1256 947 1268 981
rect 1210 941 1268 947
rect 1328 981 1386 987
rect 1328 947 1340 981
rect 1374 947 1386 981
rect 1328 941 1386 947
rect 1446 981 1504 987
rect 1446 947 1458 981
rect 1492 947 1504 981
rect 1446 941 1504 947
rect 1564 981 1622 987
rect 1564 947 1576 981
rect 1610 947 1622 981
rect 1564 941 1622 947
rect 1682 981 1740 987
rect 1682 947 1694 981
rect 1728 947 1740 981
rect 1682 941 1740 947
rect 1800 981 1858 987
rect 1800 947 1812 981
rect 1846 947 1858 981
rect 1800 941 1858 947
rect 1918 981 1976 987
rect 1918 947 1930 981
rect 1964 947 1976 981
rect 1918 941 1976 947
rect 2036 981 2094 987
rect 2036 947 2048 981
rect 2082 947 2094 981
rect 2036 941 2094 947
rect 2154 981 2212 987
rect 2154 947 2166 981
rect 2200 947 2212 981
rect 2154 941 2212 947
rect 2272 981 2330 987
rect 2272 947 2284 981
rect 2318 947 2330 981
rect 2272 941 2330 947
rect 2390 981 2448 987
rect 2390 947 2402 981
rect 2436 947 2448 981
rect 2390 941 2448 947
rect 2508 981 2566 987
rect 2508 947 2520 981
rect 2554 947 2566 981
rect 2508 941 2566 947
rect 2626 981 2684 987
rect 2626 947 2638 981
rect 2672 947 2684 981
rect 2626 941 2684 947
rect 2744 981 2802 987
rect 2744 947 2756 981
rect 2790 947 2802 981
rect 2744 941 2802 947
rect 2862 981 2920 987
rect 2862 947 2874 981
rect 2908 947 2920 981
rect 2862 941 2920 947
rect 2980 981 3038 987
rect 2980 947 2992 981
rect 3026 947 3038 981
rect 2980 941 3038 947
rect 3098 981 3156 987
rect 3098 947 3110 981
rect 3144 947 3156 981
rect 3098 941 3156 947
rect 3216 981 3274 987
rect 3216 947 3228 981
rect 3262 947 3274 981
rect 3216 941 3274 947
rect 3334 981 3392 987
rect 3334 947 3346 981
rect 3380 947 3392 981
rect 3334 941 3392 947
rect 3452 981 3510 987
rect 3452 947 3464 981
rect 3498 947 3510 981
rect 3452 941 3510 947
rect -3563 888 -3517 900
rect -3563 -888 -3557 888
rect -3523 -888 -3517 888
rect -3563 -900 -3517 -888
rect -3445 888 -3399 900
rect -3445 -888 -3439 888
rect -3405 -888 -3399 888
rect -3445 -900 -3399 -888
rect -3327 888 -3281 900
rect -3327 -888 -3321 888
rect -3287 -888 -3281 888
rect -3327 -900 -3281 -888
rect -3209 888 -3163 900
rect -3209 -888 -3203 888
rect -3169 -888 -3163 888
rect -3209 -900 -3163 -888
rect -3091 888 -3045 900
rect -3091 -888 -3085 888
rect -3051 -888 -3045 888
rect -3091 -900 -3045 -888
rect -2973 888 -2927 900
rect -2973 -888 -2967 888
rect -2933 -888 -2927 888
rect -2973 -900 -2927 -888
rect -2855 888 -2809 900
rect -2855 -888 -2849 888
rect -2815 -888 -2809 888
rect -2855 -900 -2809 -888
rect -2737 888 -2691 900
rect -2737 -888 -2731 888
rect -2697 -888 -2691 888
rect -2737 -900 -2691 -888
rect -2619 888 -2573 900
rect -2619 -888 -2613 888
rect -2579 -888 -2573 888
rect -2619 -900 -2573 -888
rect -2501 888 -2455 900
rect -2501 -888 -2495 888
rect -2461 -888 -2455 888
rect -2501 -900 -2455 -888
rect -2383 888 -2337 900
rect -2383 -888 -2377 888
rect -2343 -888 -2337 888
rect -2383 -900 -2337 -888
rect -2265 888 -2219 900
rect -2265 -888 -2259 888
rect -2225 -888 -2219 888
rect -2265 -900 -2219 -888
rect -2147 888 -2101 900
rect -2147 -888 -2141 888
rect -2107 -888 -2101 888
rect -2147 -900 -2101 -888
rect -2029 888 -1983 900
rect -2029 -888 -2023 888
rect -1989 -888 -1983 888
rect -2029 -900 -1983 -888
rect -1911 888 -1865 900
rect -1911 -888 -1905 888
rect -1871 -888 -1865 888
rect -1911 -900 -1865 -888
rect -1793 888 -1747 900
rect -1793 -888 -1787 888
rect -1753 -888 -1747 888
rect -1793 -900 -1747 -888
rect -1675 888 -1629 900
rect -1675 -888 -1669 888
rect -1635 -888 -1629 888
rect -1675 -900 -1629 -888
rect -1557 888 -1511 900
rect -1557 -888 -1551 888
rect -1517 -888 -1511 888
rect -1557 -900 -1511 -888
rect -1439 888 -1393 900
rect -1439 -888 -1433 888
rect -1399 -888 -1393 888
rect -1439 -900 -1393 -888
rect -1321 888 -1275 900
rect -1321 -888 -1315 888
rect -1281 -888 -1275 888
rect -1321 -900 -1275 -888
rect -1203 888 -1157 900
rect -1203 -888 -1197 888
rect -1163 -888 -1157 888
rect -1203 -900 -1157 -888
rect -1085 888 -1039 900
rect -1085 -888 -1079 888
rect -1045 -888 -1039 888
rect -1085 -900 -1039 -888
rect -967 888 -921 900
rect -967 -888 -961 888
rect -927 -888 -921 888
rect -967 -900 -921 -888
rect -849 888 -803 900
rect -849 -888 -843 888
rect -809 -888 -803 888
rect -849 -900 -803 -888
rect -731 888 -685 900
rect -731 -888 -725 888
rect -691 -888 -685 888
rect -731 -900 -685 -888
rect -613 888 -567 900
rect -613 -888 -607 888
rect -573 -888 -567 888
rect -613 -900 -567 -888
rect -495 888 -449 900
rect -495 -888 -489 888
rect -455 -888 -449 888
rect -495 -900 -449 -888
rect -377 888 -331 900
rect -377 -888 -371 888
rect -337 -888 -331 888
rect -377 -900 -331 -888
rect -259 888 -213 900
rect -259 -888 -253 888
rect -219 -888 -213 888
rect -259 -900 -213 -888
rect -141 888 -95 900
rect -141 -888 -135 888
rect -101 -888 -95 888
rect -141 -900 -95 -888
rect -23 888 23 900
rect -23 -888 -17 888
rect 17 -888 23 888
rect -23 -900 23 -888
rect 95 888 141 900
rect 95 -888 101 888
rect 135 -888 141 888
rect 95 -900 141 -888
rect 213 888 259 900
rect 213 -888 219 888
rect 253 -888 259 888
rect 213 -900 259 -888
rect 331 888 377 900
rect 331 -888 337 888
rect 371 -888 377 888
rect 331 -900 377 -888
rect 449 888 495 900
rect 449 -888 455 888
rect 489 -888 495 888
rect 449 -900 495 -888
rect 567 888 613 900
rect 567 -888 573 888
rect 607 -888 613 888
rect 567 -900 613 -888
rect 685 888 731 900
rect 685 -888 691 888
rect 725 -888 731 888
rect 685 -900 731 -888
rect 803 888 849 900
rect 803 -888 809 888
rect 843 -888 849 888
rect 803 -900 849 -888
rect 921 888 967 900
rect 921 -888 927 888
rect 961 -888 967 888
rect 921 -900 967 -888
rect 1039 888 1085 900
rect 1039 -888 1045 888
rect 1079 -888 1085 888
rect 1039 -900 1085 -888
rect 1157 888 1203 900
rect 1157 -888 1163 888
rect 1197 -888 1203 888
rect 1157 -900 1203 -888
rect 1275 888 1321 900
rect 1275 -888 1281 888
rect 1315 -888 1321 888
rect 1275 -900 1321 -888
rect 1393 888 1439 900
rect 1393 -888 1399 888
rect 1433 -888 1439 888
rect 1393 -900 1439 -888
rect 1511 888 1557 900
rect 1511 -888 1517 888
rect 1551 -888 1557 888
rect 1511 -900 1557 -888
rect 1629 888 1675 900
rect 1629 -888 1635 888
rect 1669 -888 1675 888
rect 1629 -900 1675 -888
rect 1747 888 1793 900
rect 1747 -888 1753 888
rect 1787 -888 1793 888
rect 1747 -900 1793 -888
rect 1865 888 1911 900
rect 1865 -888 1871 888
rect 1905 -888 1911 888
rect 1865 -900 1911 -888
rect 1983 888 2029 900
rect 1983 -888 1989 888
rect 2023 -888 2029 888
rect 1983 -900 2029 -888
rect 2101 888 2147 900
rect 2101 -888 2107 888
rect 2141 -888 2147 888
rect 2101 -900 2147 -888
rect 2219 888 2265 900
rect 2219 -888 2225 888
rect 2259 -888 2265 888
rect 2219 -900 2265 -888
rect 2337 888 2383 900
rect 2337 -888 2343 888
rect 2377 -888 2383 888
rect 2337 -900 2383 -888
rect 2455 888 2501 900
rect 2455 -888 2461 888
rect 2495 -888 2501 888
rect 2455 -900 2501 -888
rect 2573 888 2619 900
rect 2573 -888 2579 888
rect 2613 -888 2619 888
rect 2573 -900 2619 -888
rect 2691 888 2737 900
rect 2691 -888 2697 888
rect 2731 -888 2737 888
rect 2691 -900 2737 -888
rect 2809 888 2855 900
rect 2809 -888 2815 888
rect 2849 -888 2855 888
rect 2809 -900 2855 -888
rect 2927 888 2973 900
rect 2927 -888 2933 888
rect 2967 -888 2973 888
rect 2927 -900 2973 -888
rect 3045 888 3091 900
rect 3045 -888 3051 888
rect 3085 -888 3091 888
rect 3045 -900 3091 -888
rect 3163 888 3209 900
rect 3163 -888 3169 888
rect 3203 -888 3209 888
rect 3163 -900 3209 -888
rect 3281 888 3327 900
rect 3281 -888 3287 888
rect 3321 -888 3327 888
rect 3281 -900 3327 -888
rect 3399 888 3445 900
rect 3399 -888 3405 888
rect 3439 -888 3445 888
rect 3399 -900 3445 -888
rect 3517 888 3563 900
rect 3517 -888 3523 888
rect 3557 -888 3563 888
rect 3517 -900 3563 -888
rect -3510 -947 -3452 -941
rect -3510 -981 -3498 -947
rect -3464 -981 -3452 -947
rect -3510 -987 -3452 -981
rect -3392 -947 -3334 -941
rect -3392 -981 -3380 -947
rect -3346 -981 -3334 -947
rect -3392 -987 -3334 -981
rect -3274 -947 -3216 -941
rect -3274 -981 -3262 -947
rect -3228 -981 -3216 -947
rect -3274 -987 -3216 -981
rect -3156 -947 -3098 -941
rect -3156 -981 -3144 -947
rect -3110 -981 -3098 -947
rect -3156 -987 -3098 -981
rect -3038 -947 -2980 -941
rect -3038 -981 -3026 -947
rect -2992 -981 -2980 -947
rect -3038 -987 -2980 -981
rect -2920 -947 -2862 -941
rect -2920 -981 -2908 -947
rect -2874 -981 -2862 -947
rect -2920 -987 -2862 -981
rect -2802 -947 -2744 -941
rect -2802 -981 -2790 -947
rect -2756 -981 -2744 -947
rect -2802 -987 -2744 -981
rect -2684 -947 -2626 -941
rect -2684 -981 -2672 -947
rect -2638 -981 -2626 -947
rect -2684 -987 -2626 -981
rect -2566 -947 -2508 -941
rect -2566 -981 -2554 -947
rect -2520 -981 -2508 -947
rect -2566 -987 -2508 -981
rect -2448 -947 -2390 -941
rect -2448 -981 -2436 -947
rect -2402 -981 -2390 -947
rect -2448 -987 -2390 -981
rect -2330 -947 -2272 -941
rect -2330 -981 -2318 -947
rect -2284 -981 -2272 -947
rect -2330 -987 -2272 -981
rect -2212 -947 -2154 -941
rect -2212 -981 -2200 -947
rect -2166 -981 -2154 -947
rect -2212 -987 -2154 -981
rect -2094 -947 -2036 -941
rect -2094 -981 -2082 -947
rect -2048 -981 -2036 -947
rect -2094 -987 -2036 -981
rect -1976 -947 -1918 -941
rect -1976 -981 -1964 -947
rect -1930 -981 -1918 -947
rect -1976 -987 -1918 -981
rect -1858 -947 -1800 -941
rect -1858 -981 -1846 -947
rect -1812 -981 -1800 -947
rect -1858 -987 -1800 -981
rect -1740 -947 -1682 -941
rect -1740 -981 -1728 -947
rect -1694 -981 -1682 -947
rect -1740 -987 -1682 -981
rect -1622 -947 -1564 -941
rect -1622 -981 -1610 -947
rect -1576 -981 -1564 -947
rect -1622 -987 -1564 -981
rect -1504 -947 -1446 -941
rect -1504 -981 -1492 -947
rect -1458 -981 -1446 -947
rect -1504 -987 -1446 -981
rect -1386 -947 -1328 -941
rect -1386 -981 -1374 -947
rect -1340 -981 -1328 -947
rect -1386 -987 -1328 -981
rect -1268 -947 -1210 -941
rect -1268 -981 -1256 -947
rect -1222 -981 -1210 -947
rect -1268 -987 -1210 -981
rect -1150 -947 -1092 -941
rect -1150 -981 -1138 -947
rect -1104 -981 -1092 -947
rect -1150 -987 -1092 -981
rect -1032 -947 -974 -941
rect -1032 -981 -1020 -947
rect -986 -981 -974 -947
rect -1032 -987 -974 -981
rect -914 -947 -856 -941
rect -914 -981 -902 -947
rect -868 -981 -856 -947
rect -914 -987 -856 -981
rect -796 -947 -738 -941
rect -796 -981 -784 -947
rect -750 -981 -738 -947
rect -796 -987 -738 -981
rect -678 -947 -620 -941
rect -678 -981 -666 -947
rect -632 -981 -620 -947
rect -678 -987 -620 -981
rect -560 -947 -502 -941
rect -560 -981 -548 -947
rect -514 -981 -502 -947
rect -560 -987 -502 -981
rect -442 -947 -384 -941
rect -442 -981 -430 -947
rect -396 -981 -384 -947
rect -442 -987 -384 -981
rect -324 -947 -266 -941
rect -324 -981 -312 -947
rect -278 -981 -266 -947
rect -324 -987 -266 -981
rect -206 -947 -148 -941
rect -206 -981 -194 -947
rect -160 -981 -148 -947
rect -206 -987 -148 -981
rect -88 -947 -30 -941
rect -88 -981 -76 -947
rect -42 -981 -30 -947
rect -88 -987 -30 -981
rect 30 -947 88 -941
rect 30 -981 42 -947
rect 76 -981 88 -947
rect 30 -987 88 -981
rect 148 -947 206 -941
rect 148 -981 160 -947
rect 194 -981 206 -947
rect 148 -987 206 -981
rect 266 -947 324 -941
rect 266 -981 278 -947
rect 312 -981 324 -947
rect 266 -987 324 -981
rect 384 -947 442 -941
rect 384 -981 396 -947
rect 430 -981 442 -947
rect 384 -987 442 -981
rect 502 -947 560 -941
rect 502 -981 514 -947
rect 548 -981 560 -947
rect 502 -987 560 -981
rect 620 -947 678 -941
rect 620 -981 632 -947
rect 666 -981 678 -947
rect 620 -987 678 -981
rect 738 -947 796 -941
rect 738 -981 750 -947
rect 784 -981 796 -947
rect 738 -987 796 -981
rect 856 -947 914 -941
rect 856 -981 868 -947
rect 902 -981 914 -947
rect 856 -987 914 -981
rect 974 -947 1032 -941
rect 974 -981 986 -947
rect 1020 -981 1032 -947
rect 974 -987 1032 -981
rect 1092 -947 1150 -941
rect 1092 -981 1104 -947
rect 1138 -981 1150 -947
rect 1092 -987 1150 -981
rect 1210 -947 1268 -941
rect 1210 -981 1222 -947
rect 1256 -981 1268 -947
rect 1210 -987 1268 -981
rect 1328 -947 1386 -941
rect 1328 -981 1340 -947
rect 1374 -981 1386 -947
rect 1328 -987 1386 -981
rect 1446 -947 1504 -941
rect 1446 -981 1458 -947
rect 1492 -981 1504 -947
rect 1446 -987 1504 -981
rect 1564 -947 1622 -941
rect 1564 -981 1576 -947
rect 1610 -981 1622 -947
rect 1564 -987 1622 -981
rect 1682 -947 1740 -941
rect 1682 -981 1694 -947
rect 1728 -981 1740 -947
rect 1682 -987 1740 -981
rect 1800 -947 1858 -941
rect 1800 -981 1812 -947
rect 1846 -981 1858 -947
rect 1800 -987 1858 -981
rect 1918 -947 1976 -941
rect 1918 -981 1930 -947
rect 1964 -981 1976 -947
rect 1918 -987 1976 -981
rect 2036 -947 2094 -941
rect 2036 -981 2048 -947
rect 2082 -981 2094 -947
rect 2036 -987 2094 -981
rect 2154 -947 2212 -941
rect 2154 -981 2166 -947
rect 2200 -981 2212 -947
rect 2154 -987 2212 -981
rect 2272 -947 2330 -941
rect 2272 -981 2284 -947
rect 2318 -981 2330 -947
rect 2272 -987 2330 -981
rect 2390 -947 2448 -941
rect 2390 -981 2402 -947
rect 2436 -981 2448 -947
rect 2390 -987 2448 -981
rect 2508 -947 2566 -941
rect 2508 -981 2520 -947
rect 2554 -981 2566 -947
rect 2508 -987 2566 -981
rect 2626 -947 2684 -941
rect 2626 -981 2638 -947
rect 2672 -981 2684 -947
rect 2626 -987 2684 -981
rect 2744 -947 2802 -941
rect 2744 -981 2756 -947
rect 2790 -981 2802 -947
rect 2744 -987 2802 -981
rect 2862 -947 2920 -941
rect 2862 -981 2874 -947
rect 2908 -981 2920 -947
rect 2862 -987 2920 -981
rect 2980 -947 3038 -941
rect 2980 -981 2992 -947
rect 3026 -981 3038 -947
rect 2980 -987 3038 -981
rect 3098 -947 3156 -941
rect 3098 -981 3110 -947
rect 3144 -981 3156 -947
rect 3098 -987 3156 -981
rect 3216 -947 3274 -941
rect 3216 -981 3228 -947
rect 3262 -981 3274 -947
rect 3216 -987 3274 -981
rect 3334 -947 3392 -941
rect 3334 -981 3346 -947
rect 3380 -981 3392 -947
rect 3334 -987 3392 -981
rect 3452 -947 3510 -941
rect 3452 -981 3464 -947
rect 3498 -981 3510 -947
rect 3452 -987 3510 -981
<< properties >>
string FIXED_BBOX -3654 -1066 3654 1066
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 9 l 0.3 m 1 nf 60 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
